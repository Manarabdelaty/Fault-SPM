* NGSPICE file created from user_proj_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt user_proj_top clk done mc[0] mc[10] mc[11] mc[12] mc[13] mc[14] mc[15] mc[16]
+ mc[17] mc[18] mc[19] mc[1] mc[20] mc[21] mc[22] mc[23] mc[24] mc[25] mc[26] mc[27]
+ mc[28] mc[29] mc[2] mc[30] mc[31] mc[3] mc[4] mc[5] mc[6] mc[7] mc[8] mc[9] mp[0]
+ mp[10] mp[11] mp[12] mp[13] mp[14] mp[15] mp[16] mp[17] mp[18] mp[19] mp[1] mp[20]
+ mp[21] mp[22] mp[23] mp[24] mp[25] mp[26] mp[27] mp[28] mp[29] mp[2] mp[30] mp[31]
+ mp[3] mp[4] mp[5] mp[6] mp[7] mp[8] mp[9] prod[0] prod[10] prod[11] prod[12] prod[13]
+ prod[14] prod[15] prod[16] prod[17] prod[18] prod[19] prod[1] prod[20] prod[21]
+ prod[22] prod[23] prod[24] prod[25] prod[26] prod[27] prod[28] prod[29] prod[2]
+ prod[30] prod[31] prod[32] prod[33] prod[34] prod[35] prod[36] prod[37] prod[38]
+ prod[39] prod[3] prod[40] prod[41] prod[42] prod[43] prod[44] prod[45] prod[46]
+ prod[47] prod[48] prod[49] prod[4] prod[50] prod[51] prod[52] prod[53] prod[54]
+ prod[55] prod[56] prod[57] prod[58] prod[59] prod[5] prod[60] prod[61] prod[62]
+ prod[63] prod[6] prod[7] prod[8] prod[9] rst start tck tdi tdo tdo_paden_o tie[0]
+ tie[100] tie[101] tie[102] tie[103] tie[104] tie[105] tie[106] tie[107] tie[108]
+ tie[109] tie[10] tie[110] tie[111] tie[112] tie[113] tie[114] tie[115] tie[116]
+ tie[117] tie[118] tie[119] tie[11] tie[120] tie[121] tie[122] tie[123] tie[124]
+ tie[125] tie[126] tie[127] tie[128] tie[129] tie[12] tie[130] tie[131] tie[132]
+ tie[133] tie[134] tie[135] tie[136] tie[137] tie[138] tie[139] tie[13] tie[140]
+ tie[141] tie[142] tie[143] tie[144] tie[145] tie[146] tie[147] tie[148] tie[149]
+ tie[14] tie[150] tie[151] tie[152] tie[153] tie[154] tie[155] tie[156] tie[157]
+ tie[158] tie[159] tie[15] tie[160] tie[161] tie[162] tie[163] tie[164] tie[165]
+ tie[166] tie[167] tie[168] tie[169] tie[16] tie[17] tie[18] tie[19] tie[1] tie[20]
+ tie[21] tie[22] tie[23] tie[24] tie[25] tie[26] tie[27] tie[28] tie[29] tie[2] tie[30]
+ tie[31] tie[32] tie[33] tie[34] tie[35] tie[36] tie[37] tie[38] tie[39] tie[3] tie[40]
+ tie[41] tie[42] tie[43] tie[44] tie[45] tie[46] tie[47] tie[48] tie[49] tie[4] tie[50]
+ tie[51] tie[52] tie[53] tie[54] tie[55] tie[56] tie[57] tie[58] tie[59] tie[5] tie[60]
+ tie[61] tie[62] tie[63] tie[64] tie[65] tie[66] tie[67] tie[68] tie[69] tie[6] tie[70]
+ tie[71] tie[72] tie[73] tie[74] tie[75] tie[76] tie[77] tie[78] tie[79] tie[7] tie[80]
+ tie[81] tie[82] tie[83] tie[84] tie[85] tie[86] tie[87] tie[88] tie[89] tie[8] tie[90]
+ tie[91] tie[92] tie[93] tie[94] tie[95] tie[96] tie[97] tie[98] tie[99] tie[9] tms
+ trst VPWR VGND
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1505__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1506_ __dut__.__uuf__._1522_/A VGND VGND VPWR VPWR __dut__.__uuf__._1506_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_123_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2740_ rst VGND VGND VPWR VPWR __dut__._2740_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2671_ rst VGND VGND VPWR VPWR __dut__._2671_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1437_ __dut__.__uuf__._1206_/X __dut__.__uuf__._1435_/X __dut__._2299_/B
+ __dut__.__uuf__._1988_/B __dut__.__uuf__._1436_/X VGND VGND VPWR VPWR __dut__._2298_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_132_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1368_ __dut__._2329_/B VGND VGND VPWR VPWR __dut__.__uuf__._1368_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1622_ __dut__._1622_/A1 __dut__._1620_/X __dut__._1621_/X VGND VGND VPWR
+ VPWR __dut__._2871_/D sky130_fd_sc_hd__a21o_4
XFILLER_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2917__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1553_ __dut__._1553_/A __dut__._2843_/Q VGND VGND VPWR VPWR __dut__._1553_/X
+ sky130_fd_sc_hd__and2_4
Xclkbuf_4_14_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2334_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1299_ __dut__.__uuf__._1308_/A VGND VGND VPWR VPWR __dut__.__uuf__._1299_/X
+ sky130_fd_sc_hd__buf_2
Xclkbuf_opt_1_tck clkbuf_opt_2_tck/A VGND VGND VPWR VPWR clkbuf_opt_1_tck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_73_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1484_ __dut__._1374_/Y mp[2] __dut__._1483_/X VGND VGND VPWR VPWR __dut__._1484_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_133_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1415__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2105_ __dut__._2105_/A __dut__._2870_/Q VGND VGND VPWR VPWR __dut__._2105_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._3085_ __dut__._3109_/CLK __dut__._3085_/D __dut__._2533_/Y VGND VGND VPWR
+ VPWR __dut__._3085_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2036_ __dut__._2044_/A1 prod[0] __dut__._2035_/X VGND VGND VPWR VPWR __dut__._3075_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_139_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_294_ _306_/CLK _294_/D trst VGND VGND VPWR VPWR _294_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_127_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2938_ __dut__._2941_/CLK __dut__._2938_/D __dut__._2680_/Y VGND VGND VPWR
+ VPWR __dut__._2938_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2869_ __dut__._2961_/CLK __dut__._2869_/D __dut__._2749_/Y VGND VGND VPWR
+ VPWR __dut__._2869_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__290__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_psn_inst_psn_buff_206_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2202__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_32_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1995__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2340_ __dut__.__uuf__._2358_/CLK __dut__._2460_/X __dut__.__uuf__._1098_/X
+ VGND VGND VPWR VPWR prod[39] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2271_ __dut__.__uuf__._2278_/CLK __dut__._2322_/X __dut__.__uuf__._1377_/X
+ VGND VGND VPWR VPWR __dut__._2323_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_141_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1222_ __dut__._2375_/B __dut__.__uuf__._1245_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1244_/A sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2498__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1153_ __dut__.__uuf__._1161_/A VGND VGND VPWR VPWR __dut__.__uuf__._1153_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1084_ __dut__.__uuf__._1087_/A VGND VGND VPWR VPWR __dut__.__uuf__._1084_/X
+ sky130_fd_sc_hd__buf_2
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1986_ __dut__.__uuf__._1986_/A VGND VGND VPWR VPWR __dut__._2236_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2723_ rst VGND VGND VPWR VPWR __dut__._2723_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2654_ rst VGND VGND VPWR VPWR __dut__._2654_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2585_ rst VGND VGND VPWR VPWR __dut__._2585_/Y sky130_fd_sc_hd__inv_2
X__dut__._1605_ __dut__._1605_/A __dut__._2866_/Q VGND VGND VPWR VPWR __dut__._1605_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_94_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1536_ __dut__._1374_/Y mp[14] __dut__._1535_/X VGND VGND VPWR VPWR __dut__._1536_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1467_ __dut__._2509_/A __dut__._2833_/Q VGND VGND VPWR VPWR __dut__._1467_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1464__A2 mc[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1398_ __dut__._1398_/A1 __dut__._1396_/X __dut__._1397_/X VGND VGND VPWR
+ VPWR __dut__._2815_/D sky130_fd_sc_hd__a21o_4
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_12_0_tck clkbuf_3_6_0_tck/X VGND VGND VPWR VPWR clkbuf_5_25_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_42_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._3068_ clkbuf_5_5_0_tck/X __dut__._3068_/D __dut__._2550_/Y VGND VGND VPWR
+ VPWR __dut__._3068_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_128_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2019_ __dut__._2207_/A __dut__._3066_/Q VGND VGND VPWR VPWR __dut__._2019_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_139_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_277_ _194_/A _277_/D VGND VGND VPWR VPWR _277_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._2704__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_156_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1840_ __dut__._1408_/X VGND VGND VPWR VPWR __dut__.__uuf__._1844_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2404__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1771_ __dut__.__uuf__._1759_/X __dut__.__uuf__._1769_/B __dut__.__uuf__._1769_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1772_/C sky130_fd_sc_hd__o21a_4
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2614__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2323_ __dut__.__uuf__._2328_/CLK __dut__._2426_/X __dut__.__uuf__._1151_/X
+ VGND VGND VPWR VPWR prod[22] sky130_fd_sc_hd__dfrtp_4
XFILLER_145_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2254_ __dut__.__uuf__._2293_/CLK __dut__._2288_/X __dut__.__uuf__._1457_/X
+ VGND VGND VPWR VPWR __dut__._2289_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1205_ __dut__.__uuf__._1205_/A VGND VGND VPWR VPWR __dut__.__uuf__._1205_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2185_ __dut__.__uuf__._2216_/CLK __dut__._2150_/X __dut__.__uuf__._1620_/X
+ VGND VGND VPWR VPWR __dut__._2151_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1136_ __dut__.__uuf__._1132_/X __dut__.__uuf__._1129_/X prod[27]
+ prod[28] __dut__.__uuf__._1126_/X VGND VGND VPWR VPWR __dut__._2436_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1694__A2 done VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2370_ __dut__._2376_/A1 __dut__._2370_/A2 __dut__._2369_/X VGND VGND VPWR
+ VPWR __dut__._2370_/X sky130_fd_sc_hd__a21o_4
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1067_ __dut__.__uuf__._1057_/X __dut__.__uuf__._1054_/X prod[50]
+ prod[51] __dut__.__uuf__._1066_/X VGND VGND VPWR VPWR __dut__._2482_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_130_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_200_ _203_/A VGND VGND VPWR VPWR _200_/X sky130_fd_sc_hd__buf_2
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1969_ __dut__._2231_/B __dut__._2237_/B VGND VGND VPWR VPWR __dut__.__uuf__._1970_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_156_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_131_ _309_/Q VGND VGND VPWR VPWR _131_/Y sky130_fd_sc_hd__inv_2
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_tck clkbuf_3_1_0_tck/A VGND VGND VPWR VPWR clkbuf_4_3_0_tck/A sky130_fd_sc_hd__clkbuf_1
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2524__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1033__A3 prod[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_90 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2268_/A1 sky130_fd_sc_hd__buf_2
XFILLER_155_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2706_ rst VGND VGND VPWR VPWR __dut__._2706_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2637_ rst VGND VGND VPWR VPWR __dut__._2637_/Y sky130_fd_sc_hd__inv_2
X__dut__._2568_ rst VGND VGND VPWR VPWR __dut__._2568_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1519_ __dut__._2509_/A __dut__._2846_/Q VGND VGND VPWR VPWR __dut__._1519_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2499_ __dut__._2499_/A prod[58] VGND VGND VPWR VPWR __dut__._2499_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1603__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_273_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1428__A2 mc[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2609__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1513__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1823_ __dut__.__uuf__._1844_/A __dut__.__uuf__._1823_/B __dut__.__uuf__._1823_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1824_/A sky130_fd_sc_hd__or3_4
XFILLER_60_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1754_ __dut__._2151_/B __dut__._2157_/B VGND VGND VPWR VPWR __dut__.__uuf__._1755_/A
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1600__A2 mp[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1685_ __dut__.__uuf__._1678_/A __dut__.__uuf__._1683_/B __dut__.__uuf__._1661_/X
+ VGND VGND VPWR VPWR __dut__._2122_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_146_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1870_ __dut__._1870_/A1 tie[87] __dut__._1869_/X VGND VGND VPWR VPWR __dut__._2992_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3090__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2306_ __dut__.__uuf__._2334_/CLK __dut__._2392_/X __dut__.__uuf__._1199_/X
+ VGND VGND VPWR VPWR prod[5] sky130_fd_sc_hd__dfrtp_4
XFILLER_102_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2237_ __dut__.__uuf__._2240_/CLK __dut__._2254_/X __dut__.__uuf__._1532_/X
+ VGND VGND VPWR VPWR __dut__._2255_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_88_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2422_ __dut__._2422_/A1 __dut__._2422_/A2 __dut__._2421_/X VGND VGND VPWR
+ VPWR __dut__._2422_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2168_ __dut__.__uuf__._2291_/CLK __dut__._2116_/X __dut__.__uuf__._1641_/X
+ VGND VGND VPWR VPWR __dut__._2117_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2099_ VGND VGND VPWR VPWR __dut__.__uuf__._2099_/HI tie[106] sky130_fd_sc_hd__conb_1
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1119_ __dut__.__uuf__._1118_/X __dut__.__uuf__._1115_/X prod[33]
+ prod[34] __dut__.__uuf__._1111_/X VGND VGND VPWR VPWR __dut__._2448_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._2353_ __dut__._2407_/A __dut__._2353_/B VGND VGND VPWR VPWR __dut__._2353_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_141_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._2519__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1423__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2284_ __dut__._2288_/A1 __dut__._2284_/A2 __dut__._2283_/X VGND VGND VPWR
+ VPWR __dut__._2284_/X sky130_fd_sc_hd__a21o_4
XFILLER_141_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1999_ __dut__._2005_/A __dut__._3056_/Q VGND VGND VPWR VPWR __dut__._1999_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_124_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_119_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1470_ __dut__.__uuf__._1492_/A VGND VGND VPWR VPWR __dut__.__uuf__._1470_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2022_ VGND VGND VPWR VPWR __dut__.__uuf__._2022_/HI tie[29] sky130_fd_sc_hd__conb_1
XFILLER_57_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2339__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1806_ __dut__.__uuf__._1799_/A __dut__.__uuf__._1804_/B __dut__.__uuf__._1774_/X
+ VGND VGND VPWR VPWR __dut__._2166_/A2 sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1737_ __dut__.__uuf__._1737_/A VGND VGND VPWR VPWR __dut__.__uuf__._1739_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._2971_ __dut__._2985_/CLK __dut__._2971_/D __dut__._2647_/Y VGND VGND VPWR
+ VPWR __dut__._2971_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1922_ __dut__._1922_/A1 tie[113] __dut__._1921_/X VGND VGND VPWR VPWR __dut__._3018_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_147_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1668_ __dut__.__uuf__._1668_/A VGND VGND VPWR VPWR __dut__.__uuf__._1668_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_136_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1853_ __dut__._1881_/A __dut__._2983_/Q VGND VGND VPWR VPWR __dut__._1853_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2802__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1599_ __dut__.__uuf__._1602_/A VGND VGND VPWR VPWR __dut__.__uuf__._1599_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1784_ __dut__._1784_/A1 tie[44] __dut__._1783_/X VGND VGND VPWR VPWR __dut__._2949_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_121_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2405_ __dut__._2407_/A prod[11] VGND VGND VPWR VPWR __dut__._2405_/X sky130_fd_sc_hd__and2_4
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2336_ __dut__._2368_/A1 __dut__._2336_/A2 __dut__._2335_/X VGND VGND VPWR
+ VPWR __dut__._2336_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2267_ __dut__._2267_/A __dut__._2267_/B VGND VGND VPWR VPWR __dut__._2267_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_222 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2423_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_211 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2499_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_200 psn_inst_psn_buff_201/A VGND VGND VPWR VPWR __dut__._2172_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_244 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1783_/A sky130_fd_sc_hd__buf_2
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_233 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2039_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_255 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2295_/A sky130_fd_sc_hd__buf_2
X__dut__._2198_ __dut__._2200_/A1 __dut__._2198_/A2 __dut__._2197_/X VGND VGND VPWR
+ VPWR __dut__._2198_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_266 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2259_/A sky130_fd_sc_hd__buf_2
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1576__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1513__A __dut__.__uuf__._1709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_288 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2105_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_277 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1445_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_299 _236_/Y VGND VGND VPWR VPWR __dut__._2509_/A sky130_fd_sc_hd__buf_8
XANTENNA___dut__._2823__CLK __dut__._2846_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2712__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1500__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_236_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2056__A2 prod[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2159__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1522_ __dut__.__uuf__._1522_/A VGND VGND VPWR VPWR __dut__.__uuf__._1522_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1453_ __dut__.__uuf__._1440_/X __dut__.__uuf__._1435_/X __dut__._2293_/B
+ __dut__.__uuf__._1447_/X __dut__.__uuf__._1452_/X VGND VGND VPWR VPWR __dut__._2292_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_144_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2622__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1384_ __dut__.__uuf__._1383_/Y __dut__.__uuf__._1373_/X __dut__.__uuf__._1374_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1384_/X sky130_fd_sc_hd__o21a_4
XFILLER_103_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2005_ VGND VGND VPWR VPWR __dut__.__uuf__._2005_/HI tie[12] sky130_fd_sc_hd__conb_1
XFILLER_122_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2121_ __dut__._2325_/A __dut__._2121_/B VGND VGND VPWR VPWR __dut__._2121_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_25_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2052_ __dut__._2412_/A1 prod[8] __dut__._2051_/X VGND VGND VPWR VPWR __dut__._3083_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1701__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2846__CLK __dut__._2846_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2954_ __dut__._2958_/CLK __dut__._2954_/D __dut__._2664_/Y VGND VGND VPWR
+ VPWR __dut__._2954_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1905_ __dut__._2005_/A __dut__._3009_/Q VGND VGND VPWR VPWR __dut__._1905_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_147_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2885_ __dut__._3102_/CLK __dut__._2885_/D __dut__._2733_/Y VGND VGND VPWR
+ VPWR __dut__._2885_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2532__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1836_ __dut__._1836_/A1 tie[70] __dut__._1835_/X VGND VGND VPWR VPWR __dut__._2975_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_150_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1767_ __dut__._1775_/A __dut__._2940_/Q VGND VGND VPWR VPWR __dut__._1767_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_150_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1698_ __dut__._1698_/A1 tie[1] __dut__._1697_/X VGND VGND VPWR VPWR __dut__._2906_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_91_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2319_ __dut__._2325_/A __dut__._2319_/B VGND VGND VPWR VPWR __dut__._2319_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2707__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1611__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__127__A tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3001__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2617__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1505_ __dut__.__uuf__._1566_/A VGND VGND VPWR VPWR __dut__.__uuf__._1522_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_151_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2670_ rst VGND VGND VPWR VPWR __dut__._2670_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1436_ __dut__._1608_/X __dut__.__uuf__._1936_/A __dut__._2301_/B
+ __dut__.__uuf__._1423_/X VGND VGND VPWR VPWR __dut__.__uuf__._1436_/X sky130_fd_sc_hd__o22a_4
XFILLER_131_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1367_ __dut__.__uuf__._1386_/A VGND VGND VPWR VPWR __dut__.__uuf__._1367_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1621_ __dut__._2197_/A __dut__._2865_/Q VGND VGND VPWR VPWR __dut__._1621_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_132_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1552_ __dut__._1374_/Y mc[4] __dut__._1551_/X VGND VGND VPWR VPWR __dut__._1552_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1298_ __dut__.__uuf__._1283_/X __dut__.__uuf__._1297_/X __dut__._2355_/B
+ __dut__.__uuf__._1283_/X VGND VGND VPWR VPWR __dut__._2354_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1483_ __dut__._2509_/A __dut__._2837_/Q VGND VGND VPWR VPWR __dut__._1483_/X
+ sky130_fd_sc_hd__and2_4
Xclkbuf_3_6_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0___dut__.__uuf__.__clk_source__/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2104_ __dut__._2104_/A1 prod[34] __dut__._2103_/X VGND VGND VPWR VPWR __dut__._3109_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2527__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1431__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._3084_ __dut__._3109_/CLK __dut__._3084_/D __dut__._2534_/Y VGND VGND VPWR
+ VPWR __dut__._3084_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2035_ __dut__._2035_/A prod[63] VGND VGND VPWR VPWR __dut__._2035_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._3024__CLK clkbuf_5_1_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_293_ _306_/CLK _293_/D trst VGND VGND VPWR VPWR _293_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2937_ __dut__._2509_/B __dut__._2937_/D __dut__._2681_/Y VGND VGND VPWR
+ VPWR __dut__._2937_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2868_ __dut__._2961_/CLK __dut__._2868_/D __dut__._2750_/Y VGND VGND VPWR
+ VPWR __dut__._2868_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1819_ __dut__._1821_/A __dut__._2966_/Q VGND VGND VPWR VPWR __dut__._1819_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_96_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2799_ rst VGND VGND VPWR VPWR __dut__._2799_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2437__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_101_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2270_ __dut__.__uuf__._2278_/CLK __dut__._2320_/X __dut__.__uuf__._1382_/X
+ VGND VGND VPWR VPWR __dut__._2321_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_113_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1221_ __dut__.__uuf__._1221_/A VGND VGND VPWR VPWR __dut__.__uuf__._1245_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_141_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1152_ __dut__.__uuf__._1147_/X __dut__.__uuf__._1144_/X prod[22]
+ prod[23] __dut__.__uuf__._1141_/X VGND VGND VPWR VPWR __dut__._2426_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1083_ __dut__.__uuf__._1072_/X __dut__.__uuf__._1069_/X prod[45]
+ prod[46] __dut__.__uuf__._1082_/X VGND VGND VPWR VPWR __dut__._2472_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3047__CLK __dut__._3058_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1985_ __dut__.__uuf__._1985_/A __dut__.__uuf__._1985_/B __dut__.__uuf__._1985_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1986_/A sky130_fd_sc_hd__or3_4
XANTENNA___dut__._2347__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2722_ rst VGND VGND VPWR VPWR __dut__._2722_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1419_ __dut__.__uuf__._1418_/Y __dut__.__uuf__._1398_/X __dut__.__uuf__._1399_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1419_/X sky130_fd_sc_hd__o21a_4
XFILLER_144_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2653_ rst VGND VGND VPWR VPWR __dut__._2653_/Y sky130_fd_sc_hd__inv_2
X__dut__._2584_ rst VGND VGND VPWR VPWR __dut__._2584_/Y sky130_fd_sc_hd__inv_2
X__dut__._1604_ __dut__._1374_/Y mp[29] __dut__._1603_/X VGND VGND VPWR VPWR __dut__._1604_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_77_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1535_ __dut__._2509_/A __dut__._2850_/Q VGND VGND VPWR VPWR __dut__._1535_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_87_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1466_ __dut__._1466_/A1 __dut__._1464_/X __dut__._1465_/X VGND VGND VPWR
+ VPWR __dut__._2832_/D sky130_fd_sc_hd__a21o_4
XFILLER_73_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1397_ __dut__._2189_/A __dut__._2814_/Q VGND VGND VPWR VPWR __dut__._1397_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._3067_ clkbuf_5_5_0_tck/X __dut__._3067_/D __dut__._2551_/Y VGND VGND VPWR
+ VPWR __dut__._3067_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2018_ __dut__._2018_/A1 tie[161] __dut__._2017_/X VGND VGND VPWR VPWR __dut__._3066_/D
+ sky130_fd_sc_hd__a21o_4
X_276_ _194_/A _276_/D VGND VGND VPWR VPWR _276_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2720__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_149_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2167__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1770_ __dut__.__uuf__._1770_/A VGND VGND VPWR VPWR __dut__.__uuf__._1772_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_60_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2168__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2322_ __dut__.__uuf__._2328_/CLK __dut__._2424_/X __dut__.__uuf__._1153_/X
+ VGND VGND VPWR VPWR prod[21] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2630__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2253_ __dut__.__uuf__._2293_/CLK __dut__._2286_/X __dut__.__uuf__._1462_/X
+ VGND VGND VPWR VPWR __dut__._2287_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2184_ __dut__.__uuf__._2216_/CLK __dut__._2148_/X __dut__.__uuf__._1621_/X
+ VGND VGND VPWR VPWR __dut__._2149_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2340__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1204_ __dut__.__uuf__._1192_/X __dut__.__uuf__._1203_/X prod[4]
+ prod[5] __dut__.__uuf__._1200_/X VGND VGND VPWR VPWR __dut__._2390_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_101_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1135_ __dut__.__uuf__._1146_/A VGND VGND VPWR VPWR __dut__.__uuf__._1135_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1066_ __dut__.__uuf__._1126_/A VGND VGND VPWR VPWR __dut__.__uuf__._1066_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1968_ __dut__._1460_/X VGND VGND VPWR VPWR __dut__.__uuf__._1972_/B
+ sky130_fd_sc_hd__inv_2
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_130_ _130_/A VGND VGND VPWR VPWR _314_/D sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2805__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1899_ __dut__.__uuf__._1899_/A VGND VGND VPWR VPWR __dut__.__uuf__._1901_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_139_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1906__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_80 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1498_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_91 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1566_/A1 sky130_fd_sc_hd__buf_2
XFILLER_105_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2705_ rst VGND VGND VPWR VPWR __dut__._2705_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2540__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2636_ rst VGND VGND VPWR VPWR __dut__._2636_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2567_ rst VGND VGND VPWR VPWR __dut__._2567_/Y sky130_fd_sc_hd__inv_2
X__dut__._1518_ __dut__._1518_/A1 __dut__._1516_/X __dut__._1517_/X VGND VGND VPWR
+ VPWR __dut__._2845_/D sky130_fd_sc_hd__a21o_4
X__dut__._2498_ __dut__._2502_/A1 __dut__._2498_/A2 __dut__._2497_/X VGND VGND VPWR
+ VPWR __dut__._2498_/X sky130_fd_sc_hd__a21o_4
XFILLER_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1449_ __dut__._2245_/A __dut__._2827_/Q VGND VGND VPWR VPWR __dut__._1449_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2398__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2715__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_259_ _194_/A _259_/D VGND VGND VPWR VPWR _259_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_143_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2322__A1 __dut__._2332_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_266_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1193__B1 prod[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1822_ __dut__._2175_/B __dut__._2181_/B __dut__.__uuf__._1821_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1823_/C sky130_fd_sc_hd__o21ai_4
XANTENNA___dut__._2625__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1753_ __dut__._1632_/X VGND VGND VPWR VPWR __dut__.__uuf__._1757_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1684_ __dut__.__uuf__._1684_/A VGND VGND VPWR VPWR __dut__._2124_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_109_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2305_ __dut__.__uuf__._2328_/CLK __dut__._2390_/X __dut__.__uuf__._1202_/X
+ VGND VGND VPWR VPWR prod[4] sky130_fd_sc_hd__dfrtp_4
XFILLER_142_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2236_ __dut__.__uuf__._2240_/CLK __dut__._2252_/X __dut__.__uuf__._1537_/X
+ VGND VGND VPWR VPWR __dut__._2253_/B sky130_fd_sc_hd__dfrtp_4
Xclkbuf_4_11_0_tck clkbuf_3_5_0_tck/X VGND VGND VPWR VPWR clkbuf_5_23_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2421_ __dut__._2507_/A prod[19] VGND VGND VPWR VPWR __dut__._2421_/X sky130_fd_sc_hd__and2_4
XFILLER_88_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2167_ __dut__.__uuf__._2291_/CLK __dut__._2114_/X __dut__.__uuf__._1642_/X
+ VGND VGND VPWR VPWR __dut__._2115_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_141_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2098_ VGND VGND VPWR VPWR __dut__.__uuf__._2098_/HI tie[105] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1118_ __dut__.__uuf__._1162_/A VGND VGND VPWR VPWR __dut__.__uuf__._1118_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2352_ __dut__._2368_/A1 __dut__._2352_/A2 __dut__._2351_/X VGND VGND VPWR
+ VPWR __dut__._2352_/X sky130_fd_sc_hd__a21o_4
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1049_ __dut__.__uuf__._1043_/X __dut__.__uuf__._1040_/X prod[56]
+ prod[57] __dut__.__uuf__._1036_/X VGND VGND VPWR VPWR __dut__._2494_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._2283_ __dut__._2303_/A __dut__._2283_/B VGND VGND VPWR VPWR __dut__._2283_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2535__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1998_ __dut__._2004_/A1 tie[151] __dut__._1997_/X VGND VGND VPWR VPWR __dut__._3056_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_152_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2619_ rst VGND VGND VPWR VPWR __dut__._2619_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._1190__A3 prod[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._3108__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2445__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2238__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_128_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2021_ VGND VGND VPWR VPWR __dut__.__uuf__._2021_/HI tie[28] sky130_fd_sc_hd__conb_1
XFILLER_97_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1181__A3 prod[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_tck clkbuf_3_1_0_tck/A VGND VGND VPWR VPWR clkbuf_4_1_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2355__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1805_ __dut__.__uuf__._1805_/A VGND VGND VPWR VPWR __dut__._2168_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_40_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1736_ __dut__.__uuf__._1736_/A __dut__.__uuf__._1736_/B __dut__.__uuf__._1736_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1737_/A sky130_fd_sc_hd__or3_4
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2970_ __dut__._2985_/CLK __dut__._2970_/D __dut__._2648_/Y VGND VGND VPWR
+ VPWR __dut__._2970_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1921_ __dut__._2207_/A __dut__._3017_/Q VGND VGND VPWR VPWR __dut__._1921_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1667_ __dut__._2119_/B __dut__._2125_/B VGND VGND VPWR VPWR __dut__.__uuf__._1668_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_134_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1852_ __dut__._1864_/A1 tie[78] __dut__._1851_/X VGND VGND VPWR VPWR __dut__._2983_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1598_ __dut__.__uuf__._1602_/A VGND VGND VPWR VPWR __dut__.__uuf__._1598_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_136_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1783_ __dut__._1783_/A __dut__._2948_/Q VGND VGND VPWR VPWR __dut__._1783_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2219_ __dut__.__uuf__._2225_/CLK __dut__._2218_/X __dut__.__uuf__._1578_/X
+ VGND VGND VPWR VPWR __dut__._2219_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_152_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2404_ __dut__._2412_/A1 __dut__._2404_/A2 __dut__._2403_/X VGND VGND VPWR
+ VPWR __dut__._2404_/X sky130_fd_sc_hd__a21o_4
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2335_ __dut__._2407_/A __dut__._2335_/B VGND VGND VPWR VPWR __dut__._2335_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_90_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2266_ __dut__._2266_/A1 __dut__._2266_/A2 __dut__._2265_/X VGND VGND VPWR
+ VPWR __dut__._2266_/X sky130_fd_sc_hd__a21o_4
X__dut__._2197_ __dut__._2197_/A __dut__._2197_/B VGND VGND VPWR VPWR __dut__._2197_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_212 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2497_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_201 psn_inst_psn_buff_201/A VGND VGND VPWR VPWR __dut__._2222_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_245 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1781_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_223 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2081_/A sky130_fd_sc_hd__buf_2
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_234 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1881_/A sky130_fd_sc_hd__buf_2
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_267 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2257_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_289 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1817_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_256 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2293_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_278 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1553_/A sky130_fd_sc_hd__buf_2
XFILLER_145_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1576__A2 mp[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1500__A2 mp[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_131_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_229_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3080__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1704__A __dut__.__uuf__._1982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2175__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1521_ __dut__.__uuf__._1507_/X __dut__.__uuf__._1502_/X __dut__._2261_/B
+ __dut__.__uuf__._1512_/X __dut__.__uuf__._1520_/X VGND VGND VPWR VPWR __dut__._2260_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_156_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1452_ __dut__._1592_/X __dut__.__uuf__._1442_/X __dut__._2295_/B
+ __dut__.__uuf__._1448_/X VGND VGND VPWR VPWR __dut__.__uuf__._1452_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1519__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1383_ __dut__._2323_/B VGND VGND VPWR VPWR __dut__.__uuf__._1383_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_103_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2004_ VGND VGND VPWR VPWR __dut__.__uuf__._2004_/HI tie[11] sky130_fd_sc_hd__conb_1
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2120_ __dut__._2120_/A1 __dut__._2120_/A2 __dut__._2119_/X VGND VGND VPWR
+ VPWR __dut__._2120_/X sky130_fd_sc_hd__a21o_4
XFILLER_81_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2051_ __dut__._2407_/A __dut__._3082_/Q VGND VGND VPWR VPWR __dut__._2051_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_13_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1719_ __dut__.__uuf__._1719_/A VGND VGND VPWR VPWR __dut__._2136_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__._2953_ __dut__._2958_/CLK __dut__._2953_/D __dut__._2665_/Y VGND VGND VPWR
+ VPWR __dut__._2953_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1904_ __dut__._2004_/A1 tie[104] __dut__._1903_/X VGND VGND VPWR VPWR __dut__._3009_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_5_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2884_ __dut__._3102_/CLK __dut__._2884_/D __dut__._2734_/Y VGND VGND VPWR
+ VPWR __dut__._2884_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1835_ __dut__._2507_/A __dut__._2974_/Q VGND VGND VPWR VPWR __dut__._1835_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1766_ __dut__._1780_/A1 tie[35] __dut__._1765_/X VGND VGND VPWR VPWR __dut__._2940_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_150_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1697_ __dut__._2189_/A __dut__._2905_/Q VGND VGND VPWR VPWR __dut__._1697_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_3_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2318_ __dut__._2318_/A1 __dut__._2318_/A2 __dut__._2317_/X VGND VGND VPWR
+ VPWR __dut__._2318_/X sky130_fd_sc_hd__a21o_4
X__dut__._2249_ __dut__._2249_/A __dut__._2249_/B VGND VGND VPWR VPWR __dut__._2249_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2723__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2633__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1504_ __dut__.__uuf__._1486_/X __dut__.__uuf__._1502_/X __dut__._2269_/B
+ __dut__.__uuf__._1491_/X __dut__.__uuf__._1503_/X VGND VGND VPWR VPWR __dut__._2268_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1435_ __dut__.__uuf__._1480_/A VGND VGND VPWR VPWR __dut__.__uuf__._1435_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_144_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1366_ __dut__.__uuf__._1461_/A VGND VGND VPWR VPWR __dut__.__uuf__._1386_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1620_ __dut__._1374_/Y mc[6] __dut__._1619_/X VGND VGND VPWR VPWR __dut__._1620_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_132_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1551_ __dut__._2509_/A __dut__._2854_/Q VGND VGND VPWR VPWR __dut__._1551_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_0___dut__.__uuf__.__clk_source___A __dut__._2510_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1297_ __dut__.__uuf__._1291_/Y __dut__.__uuf__._1294_/X __dut__.__uuf__._1296_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1297_/X sky130_fd_sc_hd__o21a_4
XFILLER_133_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1482_ __dut__._1490_/A1 __dut__._1480_/X __dut__._1481_/X VGND VGND VPWR
+ VPWR __dut__._2836_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1476__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2813__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2808__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2103_ __dut__._2103_/A __dut__._3108_/Q VGND VGND VPWR VPWR __dut__._2103_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._3083_ __dut__._3109_/CLK __dut__._3083_/D __dut__._2535_/Y VGND VGND VPWR
+ VPWR __dut__._3083_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2034_ __dut__._2034_/A1 tie[169] __dut__._2033_/X VGND VGND VPWR VPWR __dut__._3074_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_32_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_292_ _306_/CLK _292_/D trst VGND VGND VPWR VPWR _292_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1400__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2543__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2936_ clkbuf_5_9_0_tck/X __dut__._2936_/D __dut__._2682_/Y VGND VGND VPWR
+ VPWR __dut__._2936_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2867_ __dut__._2961_/CLK __dut__._2867_/D __dut__._2751_/Y VGND VGND VPWR
+ VPWR __dut__._2867_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1818_ __dut__._1818_/A1 tie[61] __dut__._1817_/X VGND VGND VPWR VPWR __dut__._2966_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_96_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2798_ rst VGND VGND VPWR VPWR __dut__._2798_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1749_ __dut__._2189_/A __dut__._2931_/Q VGND VGND VPWR VPWR __dut__._1749_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2718__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2453__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_296_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1220_ __dut__.__uuf__._1248_/A __dut__.__uuf__._1248_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1221_/A sky130_fd_sc_hd__or2_4
XFILLER_141_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1151_ __dut__.__uuf__._1161_/A VGND VGND VPWR VPWR __dut__.__uuf__._1151_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1109__A3 prod[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1082_ __dut__.__uuf__._1126_/A VGND VGND VPWR VPWR __dut__.__uuf__._1082_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2628__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1984_ __dut__.__uuf__._1680_/A __dut__.__uuf__._1982_/B __dut__.__uuf__._1982_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1985_/C sky130_fd_sc_hd__o21a_4
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2363__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2721_ rst VGND VGND VPWR VPWR __dut__._2721_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1418_ __dut__._2309_/B VGND VGND VPWR VPWR __dut__.__uuf__._1418_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_120_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2652_ rst VGND VGND VPWR VPWR __dut__._2652_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1707__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2583_ rst VGND VGND VPWR VPWR __dut__._2583_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1349_ __dut__.__uuf__._1346_/Y __dut__.__uuf__._1347_/X __dut__.__uuf__._1348_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1349_/X sky130_fd_sc_hd__o21a_4
X__dut__._1603_ __dut__._2509_/A __dut__._2867_/Q VGND VGND VPWR VPWR __dut__._1603_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1534_ __dut__._1562_/A1 __dut__._1532_/X __dut__._1533_/X VGND VGND VPWR
+ VPWR __dut__._2849_/D sky130_fd_sc_hd__a21o_4
XFILLER_100_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1465_ __dut__._2325_/A __dut__._2821_/Q VGND VGND VPWR VPWR __dut__._1465_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_85_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1396_ __dut__._1374_/Y mc[14] __dut__._1395_/X VGND VGND VPWR VPWR __dut__._1396_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2538__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3066_ clkbuf_5_4_0_tck/X __dut__._3066_/D __dut__._2552_/Y VGND VGND VPWR
+ VPWR __dut__._3066_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2017_ __dut__._2207_/A __dut__._3065_/Q VGND VGND VPWR VPWR __dut__._2017_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_53_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_275_ _290_/CLK _275_/D VGND VGND VPWR VPWR _275_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2271__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_127_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2919_ clkbuf_5_0_0_tck/X __dut__._2919_/D __dut__._2699_/Y VGND VGND VPWR
+ VPWR __dut__._2919_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_142_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1612__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_211_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2183__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0___dut__.__uuf__.__clk_source__ clkbuf_4_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2240_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2321_ __dut__.__uuf__._2328_/CLK __dut__._2422_/X __dut__.__uuf__._1155_/X
+ VGND VGND VPWR VPWR prod[20] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2252_ __dut__.__uuf__._2293_/CLK __dut__._2284_/X __dut__.__uuf__._1468_/X
+ VGND VGND VPWR VPWR __dut__._2285_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1203_ __dut__.__uuf__._1480_/A VGND VGND VPWR VPWR __dut__.__uuf__._1203_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2183_ __dut__.__uuf__._2216_/CLK __dut__._2146_/X __dut__.__uuf__._1623_/X
+ VGND VGND VPWR VPWR __dut__._2147_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1527__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3014__CLK __dut__._3059_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1134_ __dut__.__uuf__._1134_/A VGND VGND VPWR VPWR __dut__.__uuf__._1146_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1065_ __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR __dut__.__uuf__._1126_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_28_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1967_ __dut__.__uuf__._1960_/A __dut__.__uuf__._1965_/B __dut__.__uuf__._1936_/X
+ VGND VGND VPWR VPWR __dut__._2226_/A2 sky130_fd_sc_hd__o21a_4
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1622__A __dut__.__uuf__._1628_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1898_ __dut__.__uuf__._1898_/A __dut__.__uuf__._1898_/B __dut__.__uuf__._1898_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1899_/A sky130_fd_sc_hd__or3_4
XFILLER_139_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_81 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1502_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_70 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1418_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_92 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1570_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2704_ rst VGND VGND VPWR VPWR __dut__._2704_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2635_ rst VGND VGND VPWR VPWR __dut__._2635_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2566_ rst VGND VGND VPWR VPWR __dut__._2566_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3074__D __dut__._3074_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1517_ __dut__._1557_/A __dut__._2844_/Q VGND VGND VPWR VPWR __dut__._1517_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_19_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2497_ __dut__._2497_/A prod[57] VGND VGND VPWR VPWR __dut__._2497_/X sky130_fd_sc_hd__and2_4
XFILLER_104_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1448_ __dut__._1374_/Y mc[26] __dut__._1447_/X VGND VGND VPWR VPWR __dut__._1448_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_62_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1379_ __dut__._2509_/A __dut__._2811_/Q VGND VGND VPWR VPWR __dut__._1379_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3049_ __dut__._3058_/CLK __dut__._3049_/D __dut__._2569_/Y VGND VGND VPWR
+ VPWR __dut__._3049_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_258_ _306_/CLK _258_/D VGND VGND VPWR VPWR _258_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_189_ _264_/Q _191_/B VGND VGND VPWR VPWR _263_/D sky130_fd_sc_hd__and2_4
XFILLER_143_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2731__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3037__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_161_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_259_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2167__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_49_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2086__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1821_ __dut__.__uuf__._1821_/A VGND VGND VPWR VPWR __dut__.__uuf__._1821_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1752_ __dut__.__uuf__._1745_/A __dut__.__uuf__._1750_/B __dut__.__uuf__._1720_/X
+ VGND VGND VPWR VPWR __dut__._2146_/A2 sky130_fd_sc_hd__o21a_4
XANTENNA___dut__.__uuf__._1442__A __dut__.__uuf__._1563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1683_ __dut__.__uuf__._1706_/A __dut__.__uuf__._1683_/B __dut__.__uuf__._1683_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1684_/A sky130_fd_sc_hd__or3_4
XFILLER_118_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2641__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2304_ __dut__.__uuf__._2328_/CLK __dut__._2388_/X __dut__.__uuf__._1205_/X
+ VGND VGND VPWR VPWR prod[3] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2235_ __dut__.__uuf__._2240_/CLK __dut__._2250_/X __dut__.__uuf__._1540_/X
+ VGND VGND VPWR VPWR __dut__._2251_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2420_ __dut__._2422_/A1 __dut__._2420_/A2 __dut__._2419_/X VGND VGND VPWR
+ VPWR __dut__._2420_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2166_ __dut__.__uuf__._2291_/CLK __dut__._2112_/X __dut__.__uuf__._1643_/X
+ VGND VGND VPWR VPWR __dut__._2113_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_75_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1117_ __dut__.__uuf__._1117_/A VGND VGND VPWR VPWR __dut__.__uuf__._1117_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2097_ VGND VGND VPWR VPWR __dut__.__uuf__._2097_/HI tie[104] sky130_fd_sc_hd__conb_1
XFILLER_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2351_ __dut__._2407_/A __dut__._2351_/B VGND VGND VPWR VPWR __dut__._2351_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1048_ __dut__.__uuf__._1056_/A VGND VGND VPWR VPWR __dut__.__uuf__._1048_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2282_ __dut__._2288_/A1 __dut__._2282_/A2 __dut__._2281_/X VGND VGND VPWR
+ VPWR __dut__._2282_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1997_ __dut__._2005_/A __dut__._3055_/Q VGND VGND VPWR VPWR __dut__._1997_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2551__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2618_ rst VGND VGND VPWR VPWR __dut__._2618_/Y sky130_fd_sc_hd__inv_2
X__dut__._2549_ rst VGND VGND VPWR VPWR __dut__._2549_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2726__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2445__B prod[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2461__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2020_ VGND VGND VPWR VPWR __dut__.__uuf__._2020_/HI tie[27] sky130_fd_sc_hd__conb_1
XFILLER_97_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__270__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2636__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1804_ __dut__.__uuf__._1815_/A __dut__.__uuf__._1804_/B __dut__.__uuf__._1804_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1805_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1735_ __dut__._2143_/B __dut__._2149_/B __dut__.__uuf__._1734_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1736_/C sky130_fd_sc_hd__o21ai_4
XFILLER_138_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1920_ __dut__._1920_/A1 tie[112] __dut__._1919_/X VGND VGND VPWR VPWR __dut__._3017_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_153_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1666_ __dut__._1420_/X VGND VGND VPWR VPWR __dut__.__uuf__._1670_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_147_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1851_ __dut__._1881_/A __dut__._2982_/Q VGND VGND VPWR VPWR __dut__._1851_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1597_ __dut__.__uuf__._1597_/A VGND VGND VPWR VPWR __dut__.__uuf__._1602_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2371__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1782_ __dut__._1782_/A1 tie[43] __dut__._1781_/X VGND VGND VPWR VPWR __dut__._2948_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_114_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2218_ __dut__.__uuf__._2225_/CLK __dut__._2216_/X __dut__.__uuf__._1580_/X
+ VGND VGND VPWR VPWR __dut__._2217_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_152_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2149_ VGND VGND VPWR VPWR __dut__.__uuf__._2149_/HI tie[156] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._1715__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2403_ __dut__._2407_/A prod[10] VGND VGND VPWR VPWR __dut__._2403_/X sky130_fd_sc_hd__and2_4
XFILLER_75_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2334_ __dut__._2368_/A1 __dut__._2334_/A2 __dut__._2333_/X VGND VGND VPWR
+ VPWR __dut__._2334_/X sky130_fd_sc_hd__a21o_4
XFILLER_56_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_62_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2470__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2265_ __dut__._2265_/A __dut__._2265_/B VGND VGND VPWR VPWR __dut__._2265_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2546__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_202 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2220_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2196_ __dut__._2200_/A1 __dut__._2196_/A2 __dut__._2195_/X VGND VGND VPWR
+ VPWR __dut__._2196_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_213 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2505_/A sky130_fd_sc_hd__buf_2
XFILLER_32_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_246 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1777_/A sky130_fd_sc_hd__buf_2
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_224 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2073_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_235 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1843_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_268 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2189_/A sky130_fd_sc_hd__buf_8
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_257 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2303_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_279 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1509_/A sky130_fd_sc_hd__buf_2
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_124_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2205__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_tck clkbuf_3_5_0_tck/X VGND VGND VPWR VPWR clkbuf_5_21_0_tck/A sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1520_ __dut__._1524_/X __dut__.__uuf__._1508_/X __dut__._2263_/B
+ __dut__.__uuf__._1513_/X VGND VGND VPWR VPWR __dut__.__uuf__._1520_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1451_ __dut__.__uuf__._1457_/A VGND VGND VPWR VPWR __dut__.__uuf__._1451_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1720__A __dut__.__uuf__._1828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1382_ __dut__.__uuf__._1386_/A VGND VGND VPWR VPWR __dut__.__uuf__._1382_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1535__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2003_ VGND VGND VPWR VPWR __dut__.__uuf__._2003_/HI tie[10] sky130_fd_sc_hd__conb_1
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2050_ __dut__._2412_/A1 prod[7] __dut__._2049_/X VGND VGND VPWR VPWR __dut__._3082_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA__303__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1718_ __dut__.__uuf__._1761_/A __dut__.__uuf__._1718_/B __dut__.__uuf__._1718_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1719_/A sky130_fd_sc_hd__or3_4
X__dut__._2952_ __dut__._2958_/CLK __dut__._2952_/D __dut__._2666_/Y VGND VGND VPWR
+ VPWR __dut__._2952_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1903_ __dut__._2005_/A __dut__._3008_/Q VGND VGND VPWR VPWR __dut__._1903_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1649_ __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR __dut__.__uuf__._1706_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2883_ __dut__._3102_/CLK __dut__._2883_/D __dut__._2735_/Y VGND VGND VPWR
+ VPWR __dut__._2883_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1834_ __dut__._1834_/A1 tie[69] __dut__._1833_/X VGND VGND VPWR VPWR __dut__._2974_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2892__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1765_ __dut__._1775_/A __dut__._2939_/Q VGND VGND VPWR VPWR __dut__._1765_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1696_ __dut__._1696_/A1 tie[0] __dut__._1695_/X VGND VGND VPWR VPWR __dut__._2905_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2228__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_91_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2317_ __dut__._2325_/A __dut__._2317_/B VGND VGND VPWR VPWR __dut__._2317_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_17_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2248_ __dut__._2250_/A1 __dut__._2248_/A2 __dut__._2247_/X VGND VGND VPWR
+ VPWR __dut__._2248_/X sky130_fd_sc_hd__a21o_4
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2179_ __dut__._2189_/A __dut__._2179_/B VGND VGND VPWR VPWR __dut__._2179_/X
+ sky130_fd_sc_hd__and2_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_241_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1503_ __dut__._1540_/X __dut__.__uuf__._1487_/X __dut__._2271_/B
+ __dut__.__uuf__._1492_/X VGND VGND VPWR VPWR __dut__.__uuf__._1503_/X sky130_fd_sc_hd__o22a_4
XFILLER_116_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1434_ __dut__.__uuf__._1434_/A VGND VGND VPWR VPWR __dut__.__uuf__._1434_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_117_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1365_ __dut__.__uuf__._1603_/A VGND VGND VPWR VPWR __dut__.__uuf__._1461_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_89_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1550_ __dut__._1562_/A1 __dut__._1548_/X __dut__._1549_/X VGND VGND VPWR
+ VPWR __dut__._2853_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1296_ __dut__.__uuf__._1322_/A VGND VGND VPWR VPWR __dut__.__uuf__._1296_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1476__A2 mp[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1481_ __dut__._2281_/A __dut__._2835_/Q VGND VGND VPWR VPWR __dut__._1481_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2102_ __dut__._2102_/A1 prod[33] __dut__._2101_/X VGND VGND VPWR VPWR __dut__._3108_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._3082_ __dut__._3093_/CLK __dut__._3082_/D __dut__._2536_/Y VGND VGND VPWR
+ VPWR __dut__._3082_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2033_ __dut__._2207_/A __dut__._3073_/Q VGND VGND VPWR VPWR __dut__._2033_/X
+ sky130_fd_sc_hd__and2_4
X_291_ _306_/CLK _291_/D trst VGND VGND VPWR VPWR _291_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_25_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1400__A2 mc[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2935_ clkbuf_5_9_0_tck/X __dut__._2935_/D __dut__._2683_/Y VGND VGND VPWR
+ VPWR __dut__._2935_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2866_ __dut__._2961_/CLK __dut__._2866_/D __dut__._2752_/Y VGND VGND VPWR
+ VPWR __dut__._2866_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1817_ __dut__._1817_/A __dut__._2965_/Q VGND VGND VPWR VPWR __dut__._1817_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._3070__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2797_ rst VGND VGND VPWR VPWR __dut__._2797_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1748_ __dut__._1942_/A1 tie[26] __dut__._1747_/X VGND VGND VPWR VPWR __dut__._2931_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__296__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1679_ __dut__._1891_/A __dut__._2896_/Q VGND VGND VPWR VPWR __dut__._1679_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1903__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2734__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2453__B prod[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_289_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_191_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1150_ __dut__.__uuf__._1208_/A VGND VGND VPWR VPWR __dut__.__uuf__._1161_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_141_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1081_ __dut__.__uuf__._1087_/A VGND VGND VPWR VPWR __dut__.__uuf__._1081_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1983_ __dut__.__uuf__._1983_/A VGND VGND VPWR VPWR __dut__.__uuf__._1985_/B
+ sky130_fd_sc_hd__inv_2
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2644__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3093__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2720_ rst VGND VGND VPWR VPWR __dut__._2720_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2651_ rst VGND VGND VPWR VPWR __dut__._2651_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1417_ __dut__.__uuf__._1434_/A VGND VGND VPWR VPWR __dut__.__uuf__._1417_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1602_ __dut__._1780_/A1 __dut__._1600_/X __dut__._1601_/X VGND VGND VPWR
+ VPWR __dut__._2866_/D sky130_fd_sc_hd__a21o_4
XFILLER_144_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2582_ rst VGND VGND VPWR VPWR __dut__._2582_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1348_ __dut__.__uuf__._1399_/A VGND VGND VPWR VPWR __dut__.__uuf__._1348_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1533_ __dut__._1557_/A __dut__._2848_/Q VGND VGND VPWR VPWR __dut__._1533_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1279_ __dut__.__uuf__._1271_/X __dut__.__uuf__._1278_/X __dut__._2361_/B
+ __dut__.__uuf__._1271_/X VGND VGND VPWR VPWR __dut__._2360_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1464_ __dut__._1374_/Y mc[2] __dut__._1463_/X VGND VGND VPWR VPWR __dut__._1464_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_37_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1723__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1395_ __dut__._2509_/A __dut__._2815_/Q VGND VGND VPWR VPWR __dut__._1395_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3065_ clkbuf_5_4_0_tck/X __dut__._3065_/D __dut__._2553_/Y VGND VGND VPWR
+ VPWR __dut__._3065_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2016_ __dut__._2016_/A1 tie[160] __dut__._2015_/X VGND VGND VPWR VPWR __dut__._3065_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2554__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_274_ _274_/CLK _274_/D VGND VGND VPWR VPWR _274_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2918_ clkbuf_5_0_0_tck/X __dut__._2918_/D __dut__._2700_/Y VGND VGND VPWR
+ VPWR __dut__._2918_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2849_ __dut__._2860_/CLK __dut__._2849_/D __dut__._2769_/Y VGND VGND VPWR
+ VPWR __dut__._2849_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1688__A2 prod[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2729__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1612__A2 mp[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1376__A1 mc[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2320_ __dut__.__uuf__._2328_/CLK __dut__._2420_/X __dut__.__uuf__._1158_/X
+ VGND VGND VPWR VPWR prod[19] sky130_fd_sc_hd__dfrtp_4
XFILLER_114_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2251_ __dut__.__uuf__._2251_/CLK __dut__._2282_/X __dut__.__uuf__._1473_/X
+ VGND VGND VPWR VPWR __dut__._2283_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1202_ __dut__.__uuf__._1205_/A VGND VGND VPWR VPWR __dut__.__uuf__._1202_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_102_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2182_ __dut__.__uuf__._2216_/CLK __dut__._2144_/X __dut__.__uuf__._1624_/X
+ VGND VGND VPWR VPWR __dut__._2145_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1133_ __dut__.__uuf__._1132_/X __dut__.__uuf__._1129_/X prod[28]
+ prod[29] __dut__.__uuf__._1126_/X VGND VGND VPWR VPWR __dut__._2438_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_101_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1064_ __dut__.__uuf__._1071_/A VGND VGND VPWR VPWR __dut__.__uuf__._1064_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1543__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2639__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1966_ __dut__.__uuf__._1966_/A VGND VGND VPWR VPWR __dut__._2228_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1897_ __dut__._2203_/B __dut__._2209_/B __dut__.__uuf__._1896_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1898_/C sky130_fd_sc_hd__o21ai_4
XFILLER_137_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2703_ rst VGND VGND VPWR VPWR __dut__._2703_/Y sky130_fd_sc_hd__inv_2
Xpsn_inst_psn_buff_82 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1506_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_71 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1430_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_60 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1474_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_151_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_93 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2294_/A1 sky130_fd_sc_hd__buf_2
XFILLER_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2634_ rst VGND VGND VPWR VPWR __dut__._2634_/Y sky130_fd_sc_hd__inv_2
X__dut__._2565_ rst VGND VGND VPWR VPWR __dut__._2565_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_10_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2353_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA_psn_inst_psn_buff_92_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1516_ __dut__._1374_/Y mp[9] __dut__._1515_/X VGND VGND VPWR VPWR __dut__._1516_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_19_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2549__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2496_ __dut__._2502_/A1 __dut__._2496_/A2 __dut__._2495_/X VGND VGND VPWR
+ VPWR __dut__._2496_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1453__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1447_ __dut__._2509_/A __dut__._2828_/Q VGND VGND VPWR VPWR __dut__._1447_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_27_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1378_ __dut__._2288_/A1 __dut__._1376_/X __dut__._1377_/X VGND VGND VPWR
+ VPWR __dut__._2810_/D sky130_fd_sc_hd__a21o_4
X__dut__._3048_ __dut__._3058_/CLK __dut__._3048_/D __dut__._2570_/Y VGND VGND VPWR
+ VPWR __dut__._3048_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_257_ _306_/CLK _257_/D VGND VGND VPWR VPWR _258_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_155_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_188_ _265_/Q _191_/B VGND VGND VPWR VPWR _264_/D sky130_fd_sc_hd__and2_4
XFILLER_89_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2459__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_154_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1820_ __dut__._2175_/B __dut__._2181_/B VGND VGND VPWR VPWR __dut__.__uuf__._1821_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_33_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1751_ __dut__.__uuf__._1751_/A VGND VGND VPWR VPWR __dut__._2148_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1682_ __dut__.__uuf__._1261_/X __dut__.__uuf__._1680_/B __dut__.__uuf__._1680_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1683_/C sky130_fd_sc_hd__o21a_4
XFILLER_119_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2303_ __dut__.__uuf__._2303_/CLK __dut__._2386_/X __dut__.__uuf__._1209_/X
+ VGND VGND VPWR VPWR prod[2] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2234_ __dut__.__uuf__._2240_/CLK __dut__._2248_/X __dut__.__uuf__._1543_/X
+ VGND VGND VPWR VPWR __dut__._2249_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2165_ __dut__.__uuf__._2291_/CLK __dut__._2110_/X __dut__.__uuf__._1644_/X
+ VGND VGND VPWR VPWR __dut__._2111_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1116_ __dut__.__uuf__._1103_/X __dut__.__uuf__._1115_/X prod[34]
+ prod[35] __dut__.__uuf__._1111_/X VGND VGND VPWR VPWR __dut__._2450_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._2096_ VGND VGND VPWR VPWR __dut__.__uuf__._2096_/HI tie[103] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2369__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2350_ __dut__._2368_/A1 __dut__._2350_/A2 __dut__._2349_/X VGND VGND VPWR
+ VPWR __dut__._2350_/X sky130_fd_sc_hd__a21o_4
XFILLER_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1047_ __dut__.__uuf__._1043_/X __dut__.__uuf__._1040_/X prod[57]
+ prod[58] __dut__.__uuf__._1036_/X VGND VGND VPWR VPWR __dut__._2496_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._2281_ __dut__._2281_/A __dut__._2281_/B VGND VGND VPWR VPWR __dut__._2281_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2849__CLK __dut__._2860_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1588__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1949_ __dut__._2223_/B __dut__._2229_/B VGND VGND VPWR VPWR __dut__.__uuf__._1950_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1996_ __dut__._2004_/A1 tie[150] __dut__._1995_/X VGND VGND VPWR VPWR __dut__._3055_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_152_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2617_ rst VGND VGND VPWR VPWR __dut__._2617_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1512__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2548_ rst VGND VGND VPWR VPWR __dut__._2548_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_5_31_0_tck clkbuf_5_31_0_tck/A VGND VGND VPWR VPWR __dut__._3058_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2479_ __dut__._2491_/A prod[48] VGND VGND VPWR VPWR __dut__._2479_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1911__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_309_ _315_/CLK _309_/D trst VGND VGND VPWR VPWR _309_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2742__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_271_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2189__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1803_ __dut__.__uuf__._1759_/X __dut__.__uuf__._1801_/B __dut__.__uuf__._1801_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1804_/C sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1734_ __dut__.__uuf__._1734_/A VGND VGND VPWR VPWR __dut__.__uuf__._1734_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_138_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2652__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1665_ __dut__._2115_/B __dut__.__uuf__._1663_/X __dut__._2114_/A2
+ VGND VGND VPWR VPWR __dut__._2116_/A2 sky130_fd_sc_hd__a21boi_4
X__dut__._1850_ __dut__._1864_/A1 tie[77] __dut__._1849_/X VGND VGND VPWR VPWR __dut__._2982_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1596_ __dut__.__uuf__._1596_/A VGND VGND VPWR VPWR __dut__.__uuf__._1596_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_134_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1781_ __dut__._1781_/A __dut__._2947_/Q VGND VGND VPWR VPWR __dut__._1781_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_136_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2217_ __dut__.__uuf__._2225_/CLK __dut__._2214_/X __dut__.__uuf__._1581_/X
+ VGND VGND VPWR VPWR __dut__._2215_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_76_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2148_ VGND VGND VPWR VPWR __dut__.__uuf__._2148_/HI tie[155] sky130_fd_sc_hd__conb_1
XANTENNA___dut__.__uuf__._1628__A __dut__.__uuf__._1628_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2402_ __dut__._2412_/A1 __dut__._2402_/A2 __dut__._2401_/X VGND VGND VPWR
+ VPWR __dut__._2402_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2099__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2333_ __dut__._2407_/A __dut__._2333_/B VGND VGND VPWR VPWR __dut__._2333_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._2079_ VGND VGND VPWR VPWR __dut__.__uuf__._2079_/HI tie[86] sky130_fd_sc_hd__conb_1
XFILLER_28_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1731__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2264_ __dut__._2264_/A1 __dut__._2264_/A2 __dut__._2263_/X VGND VGND VPWR
+ VPWR __dut__._2264_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_203 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1990_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._3027__CLK clkbuf_5_1_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2195_ __dut__._2197_/A __dut__._2195_/B VGND VGND VPWR VPWR __dut__._2195_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_101_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_236 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1829_/A sky130_fd_sc_hd__buf_2
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_225 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2071_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_214 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2457_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_247 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1779_/A sky130_fd_sc_hd__buf_2
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0___dut__.__uuf__.__clk_source__ clkbuf_4_9_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2303_/CLK sky130_fd_sc_hd__clkbuf_1
Xpsn_inst_psn_buff_269 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2255_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_258 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1573_/A sky130_fd_sc_hd__buf_2
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2562__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1979_ __dut__._2005_/A __dut__._3046_/Q VGND VGND VPWR VPWR __dut__._1979_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_125_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0___dut__.__uuf__.__clk_source__ clkbuf_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR clkbuf_2_3_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_94_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2737__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__157__A tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_117_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1972__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1450_ __dut__.__uuf__._1440_/X __dut__.__uuf__._1435_/X __dut__._2295_/B
+ __dut__.__uuf__._1447_/X __dut__.__uuf__._1449_/X VGND VGND VPWR VPWR __dut__._2294_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_143_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1381_ __dut__.__uuf__._1378_/X __dut__.__uuf__._1380_/X __dut__._2323_/B
+ __dut__.__uuf__._1378_/X VGND VGND VPWR VPWR __dut__._2322_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2002_ VGND VGND VPWR VPWR __dut__.__uuf__._2002_/HI tie[9] sky130_fd_sc_hd__conb_1
XFILLER_73_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2647__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1551__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1717_ __dut__.__uuf__._1704_/X __dut__.__uuf__._1715_/B __dut__.__uuf__._1715_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1718_/C sky130_fd_sc_hd__o21a_4
X__dut__._2951_ __dut__._2958_/CLK __dut__._2951_/D __dut__._2667_/Y VGND VGND VPWR
+ VPWR __dut__._2951_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1902_ __dut__._2004_/A1 tie[103] __dut__._1901_/X VGND VGND VPWR VPWR __dut__._3008_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2882_ __dut__._3102_/CLK __dut__._2882_/D __dut__._2736_/Y VGND VGND VPWR
+ VPWR __dut__._2882_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1648_ __dut__.__uuf__._1648_/A VGND VGND VPWR VPWR done sky130_fd_sc_hd__buf_2
X__dut__._1833_ __dut__._2507_/A __dut__._2973_/Q VGND VGND VPWR VPWR __dut__._1833_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_107_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1579_ __dut__.__uuf__._1597_/A VGND VGND VPWR VPWR __dut__.__uuf__._1584_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1764_ __dut__._1780_/A1 tie[34] __dut__._1763_/X VGND VGND VPWR VPWR __dut__._2939_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1695_ __dut__._2189_/A __dut__._2904_/Q VGND VGND VPWR VPWR __dut__._1695_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_103_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2557__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2316_ __dut__._2318_/A1 __dut__._2316_/A2 __dut__._2315_/X VGND VGND VPWR
+ VPWR __dut__._2316_/X sky130_fd_sc_hd__a21o_4
X__dut__._2247_ __dut__._2247_/A __dut__._2247_/B VGND VGND VPWR VPWR __dut__._2247_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_32_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1461__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2178_ __dut__._2184_/A1 __dut__._2178_/A2 __dut__._2177_/X VGND VGND VPWR
+ VPWR __dut__._2178_/X sky130_fd_sc_hd__a21o_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2467__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_234_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1502_ __dut__.__uuf__._1563_/A VGND VGND VPWR VPWR __dut__.__uuf__._1502_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1433_ __dut__.__uuf__._1255_/X __dut__.__uuf__._1432_/X __dut__._2301_/B
+ __dut__.__uuf__._1255_/X VGND VGND VPWR VPWR __dut__._2300_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1364_ __dut__.__uuf__._1352_/X __dut__.__uuf__._1362_/X __dut__._2329_/B
+ __dut__.__uuf__._1363_/X VGND VGND VPWR VPWR __dut__._2328_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1295_ __dut__.__uuf__._1399_/A VGND VGND VPWR VPWR __dut__.__uuf__._1322_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2122__A1 __dut__._2332_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1480_ __dut__._1374_/Y mp[1] __dut__._1479_/X VGND VGND VPWR VPWR __dut__._1480_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_85_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2377__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3081_ __dut__._3093_/CLK __dut__._3081_/D __dut__._2537_/Y VGND VGND VPWR
+ VPWR __dut__._3081_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2101_ __dut__._2507_/A __dut__._3107_/Q VGND VGND VPWR VPWR __dut__._2101_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2032_ __dut__._2032_/A1 tie[168] __dut__._2031_/X VGND VGND VPWR VPWR __dut__._3073_/D
+ sky130_fd_sc_hd__a21o_4
X_290_ _290_/CLK _290_/D VGND VGND VPWR VPWR _290_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__283__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_18_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2934_ clkbuf_5_9_0_tck/X __dut__._2934_/D __dut__._2684_/Y VGND VGND VPWR
+ VPWR __dut__._2934_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2865_ clkbuf_5_3_0_tck/X __dut__._2865_/D __dut__._2753_/Y VGND VGND VPWR
+ VPWR __dut__._2865_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1816_ __dut__._1816_/A1 tie[60] __dut__._1815_/X VGND VGND VPWR VPWR __dut__._2965_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2796_ rst VGND VGND VPWR VPWR __dut__._2796_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1747_ __dut__._2189_/A __dut__._2930_/Q VGND VGND VPWR VPWR __dut__._1747_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_67_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1678_ __dut__._2502_/A1 prod[56] __dut__._1677_/X VGND VGND VPWR VPWR __dut__._2896_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2750__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2352__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1080_ __dut__.__uuf__._1072_/X __dut__.__uuf__._1069_/X prod[46]
+ prod[47] __dut__.__uuf__._1066_/X VGND VGND VPWR VPWR __dut__._2474_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_67_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1982_ __dut__.__uuf__._1982_/A __dut__.__uuf__._1982_/B __dut__.__uuf__._1982_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1983_/A sky130_fd_sc_hd__or3_4
XFILLER_36_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2882__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2660__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2650_ rst VGND VGND VPWR VPWR __dut__._2650_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1416_ __dut__.__uuf__._1461_/A VGND VGND VPWR VPWR __dut__.__uuf__._1434_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_132_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1347_ __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR __dut__.__uuf__._1347_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1601_ __dut__._1601_/A __dut__._2864_/Q VGND VGND VPWR VPWR __dut__._1601_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_120_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2581_ rst VGND VGND VPWR VPWR __dut__._2581_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1532_ __dut__._1374_/Y mp[13] __dut__._1531_/X VGND VGND VPWR VPWR __dut__._1532_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1278_ __dut__.__uuf__._1277_/Y __dut__.__uuf__._1985_/A __dut__.__uuf__._1268_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1278_/X sky130_fd_sc_hd__o21a_4
XFILLER_74_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1463_ __dut__._2509_/A __dut__._2832_/Q VGND VGND VPWR VPWR __dut__._1463_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_37_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1394_ __dut__._1394_/A1 __dut__._1392_/X __dut__._1393_/X VGND VGND VPWR
+ VPWR __dut__._2814_/D sky130_fd_sc_hd__a21o_4
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3064_ clkbuf_5_4_0_tck/X __dut__._3064_/D __dut__._2554_/Y VGND VGND VPWR
+ VPWR __dut__._3064_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2015_ __dut__._2207_/A __dut__._3064_/Q VGND VGND VPWR VPWR __dut__._2015_/X
+ sky130_fd_sc_hd__and2_4
X_273_ _274_/CLK _273_/D VGND VGND VPWR VPWR _273_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2570__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2917_ clkbuf_5_9_0_tck/X __dut__._2917_/D __dut__._2701_/Y VGND VGND VPWR
+ VPWR __dut__._2917_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._2334__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2848_ __dut__._2860_/CLK __dut__._2848_/D __dut__._2770_/Y VGND VGND VPWR
+ VPWR __dut__._2848_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2779_ rst VGND VGND VPWR VPWR __dut__._2779_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2745__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1376__A2 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1196__B1 prod[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2250_ __dut__.__uuf__._2251_/CLK __dut__._2280_/X __dut__.__uuf__._1476_/X
+ VGND VGND VPWR VPWR __dut__._2281_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_142_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1201_ __dut__.__uuf__._1192_/X __dut__.__uuf__._1189_/X prod[5]
+ prod[6] __dut__.__uuf__._1200_/X VGND VGND VPWR VPWR __dut__._2392_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_102_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2181_ __dut__.__uuf__._2216_/CLK __dut__._2142_/X __dut__.__uuf__._1625_/X
+ VGND VGND VPWR VPWR __dut__._2143_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1132_ __dut__.__uuf__._1162_/A VGND VGND VPWR VPWR __dut__.__uuf__._1132_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1063_ __dut__.__uuf__._1057_/X __dut__.__uuf__._1054_/X prod[51]
+ prod[52] __dut__.__uuf__._1051_/X VGND VGND VPWR VPWR __dut__._2484_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_83_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2655__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1965_ __dut__.__uuf__._1975_/A __dut__.__uuf__._1965_/B __dut__.__uuf__._1965_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1966_/A sky130_fd_sc_hd__or3_4
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3060__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1896_ __dut__.__uuf__._1896_/A VGND VGND VPWR VPWR __dut__.__uuf__._1896_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_83 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1514_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2702_ rst VGND VGND VPWR VPWR __dut__._2702_/Y sky130_fd_sc_hd__inv_2
Xpsn_inst_psn_buff_72 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2250_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_61 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1478_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2190__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_50 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2112_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_151_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_94 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2292_/A1 sky130_fd_sc_hd__buf_2
XFILLER_132_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2633_ rst VGND VGND VPWR VPWR __dut__._2633_/Y sky130_fd_sc_hd__inv_2
X__dut__._2564_ rst VGND VGND VPWR VPWR __dut__._2564_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0___dut__.__uuf__.__clk_source__ clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_5_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_psn_inst_psn_buff_85_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1515_ __dut__._2509_/A __dut__._2845_/Q VGND VGND VPWR VPWR __dut__._1515_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2495_ __dut__._2497_/A prod[56] VGND VGND VPWR VPWR __dut__._2495_/X sky130_fd_sc_hd__and2_4
XFILLER_74_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1446_ __dut__._1446_/A1 __dut__._1444_/X __dut__._1445_/X VGND VGND VPWR
+ VPWR __dut__._2827_/D sky130_fd_sc_hd__a21o_4
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1377_ tdi __dut__._2407_/A VGND VGND VPWR VPWR __dut__._1377_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2565__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3047_ __dut__._3058_/CLK __dut__._3047_/D __dut__._2571_/Y VGND VGND VPWR
+ VPWR __dut__._3047_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_6_0___dut__.__uuf__.__clk_source___A clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_256_ _306_/CLK _256_/D VGND VGND VPWR VPWR _257_/D sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1909__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_187_ _266_/Q _187_/B VGND VGND VPWR VPWR _265_/D sky130_fd_sc_hd__or2_4
XFILLER_155_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1193__A3 prod[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_147_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3083__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1750_ __dut__.__uuf__._1761_/A __dut__.__uuf__._1750_/B __dut__.__uuf__._1750_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1751_/A sky130_fd_sc_hd__or3_4
XANTENNA___dut__._2475__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1681_ __dut__.__uuf__._1681_/A VGND VGND VPWR VPWR __dut__.__uuf__._1683_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_146_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2302_ __dut__.__uuf__._2303_/CLK __dut__._2384_/X __dut__.__uuf__._1211_/X
+ VGND VGND VPWR VPWR prod[1] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2233_ __dut__.__uuf__._2240_/CLK __dut__._2246_/X __dut__.__uuf__._1548_/X
+ VGND VGND VPWR VPWR __dut__._2247_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_114_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2164_ __dut__.__uuf__._2291_/CLK __dut__._2108_/X __dut__.__uuf__._1645_/X
+ VGND VGND VPWR VPWR __dut__._2109_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1115_ __dut__.__uuf__._1173_/A VGND VGND VPWR VPWR __dut__.__uuf__._1115_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2095_ VGND VGND VPWR VPWR __dut__.__uuf__._2095_/HI tie[102] sky130_fd_sc_hd__conb_1
XFILLER_68_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1046_ __dut__.__uuf__._1056_/A VGND VGND VPWR VPWR __dut__.__uuf__._1046_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2280_ __dut__._2288_/A1 __dut__._2280_/A2 __dut__._2279_/X VGND VGND VPWR
+ VPWR __dut__._2280_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1588__A2 mp[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1948_ __dut__._1452_/X VGND VGND VPWR VPWR __dut__.__uuf__._1952_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_156_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1879_ __dut__.__uuf__._1867_/X __dut__.__uuf__._1877_/B __dut__.__uuf__._1877_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1880_/C sky130_fd_sc_hd__o21a_4
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1729__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1995_ __dut__._2005_/A __dut__._3054_/Q VGND VGND VPWR VPWR __dut__._1995_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_137_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1512__A2 mp[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2616_ rst VGND VGND VPWR VPWR __dut__._2616_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2547_ rst VGND VGND VPWR VPWR __dut__._2547_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2478_ __dut__._2488_/A1 __dut__._2478_/A2 __dut__._2477_/X VGND VGND VPWR
+ VPWR __dut__._2478_/X sky130_fd_sc_hd__a21o_4
XFILLER_75_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1429_ __dut__._1429_/A __dut__._2822_/Q VGND VGND VPWR VPWR __dut__._1429_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_308_ _315_/CLK _308_/D trst VGND VGND VPWR VPWR _308_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_156_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_239_ _239_/A _302_/Q _239_/C VGND VGND VPWR VPWR _251_/D sky130_fd_sc_hd__or3_4
XFILLER_115_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_264_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1374__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1802_ __dut__.__uuf__._1802_/A VGND VGND VPWR VPWR __dut__.__uuf__._1804_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_139_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1733_ __dut__._2143_/B __dut__._2149_/B VGND VGND VPWR VPWR __dut__.__uuf__._1734_/A
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1664_ __dut__._2115_/B __dut__.__uuf__._1663_/X __dut__.__uuf__._1936_/A
+ VGND VGND VPWR VPWR __dut__._2114_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1595_ __dut__.__uuf__._1596_/A VGND VGND VPWR VPWR __dut__.__uuf__._1595_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_134_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1780_ __dut__._1780_/A1 tie[42] __dut__._1779_/X VGND VGND VPWR VPWR __dut__._2947_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_88_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2216_ __dut__.__uuf__._2216_/CLK __dut__._2212_/X __dut__.__uuf__._1582_/X
+ VGND VGND VPWR VPWR __dut__._2213_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2147_ VGND VGND VPWR VPWR __dut__.__uuf__._2147_/HI tie[154] sky130_fd_sc_hd__conb_1
XFILLER_76_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2401_ __dut__._2407_/A prod[9] VGND VGND VPWR VPWR __dut__._2401_/X sky130_fd_sc_hd__and2_4
XFILLER_29_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2332_ __dut__._2332_/A1 __dut__._2332_/A2 __dut__._2331_/X VGND VGND VPWR
+ VPWR __dut__._2332_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2078_ VGND VGND VPWR VPWR __dut__.__uuf__._2078_/HI tie[85] sky130_fd_sc_hd__conb_1
XFILLER_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2263_ __dut__._2263_/A __dut__._2263_/B VGND VGND VPWR VPWR __dut__._2263_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1029_ __dut__.__uuf__._1603_/A VGND VGND VPWR VPWR __dut__.__uuf__._1992_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_204 _244_/X VGND VGND VPWR VPWR __dut__._2507_/A sky130_fd_sc_hd__buf_8
X__dut__._2194_ __dut__._2200_/A1 __dut__._2194_/A2 __dut__._2193_/X VGND VGND VPWR
+ VPWR __dut__._2194_/X sky130_fd_sc_hd__a21o_4
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_237 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1825_/A sky130_fd_sc_hd__buf_2
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_226 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2419_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_215 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2407_/A sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_248 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1775_/A sky130_fd_sc_hd__buf_2
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_259 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1569_/A sky130_fd_sc_hd__buf_2
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1459__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1978_ __dut__._2004_/A1 tie[141] __dut__._1977_/X VGND VGND VPWR VPWR __dut__._3046_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1819__A __dut__._1400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2753__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2903__D __dut__._2903_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1380_ __dut__.__uuf__._1379_/Y __dut__.__uuf__._1373_/X __dut__.__uuf__._1374_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1380_/X sky130_fd_sc_hd__o21a_4
XFILLER_144_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2839__CLK __dut__._2846_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2001_ VGND VGND VPWR VPWR __dut__.__uuf__._2001_/HI tie[8] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._1488__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1464__A __dut__.__uuf__._1464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1660__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1412__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2663__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1716_ __dut__.__uuf__._1716_/A VGND VGND VPWR VPWR __dut__.__uuf__._1718_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._2950_ __dut__._2958_/CLK __dut__._2950_/D __dut__._2668_/Y VGND VGND VPWR
+ VPWR __dut__._2950_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1901_ __dut__._2005_/A __dut__._3007_/Q VGND VGND VPWR VPWR __dut__._1901_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2881_ __dut__._3106_/CLK __dut__._2881_/D __dut__._2737_/Y VGND VGND VPWR
+ VPWR __dut__._2881_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1647_ __dut__.__uuf__._1989_/A __dut__._2109_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1648_/A sky130_fd_sc_hd__and2_4
XFILLER_135_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_30_0_tck clkbuf_5_31_0_tck/A VGND VGND VPWR VPWR _274_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__._1832_ __dut__._1832_/A1 tie[68] __dut__._1831_/X VGND VGND VPWR VPWR __dut__._2973_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1578_ __dut__.__uuf__._1578_/A VGND VGND VPWR VPWR __dut__.__uuf__._1578_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1763_ __dut__._1775_/A __dut__._2938_/Q VGND VGND VPWR VPWR __dut__._1763_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1694_ __dut__._2376_/A1 done __dut__._1693_/X VGND VGND VPWR VPWR __dut__._2904_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_130_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2315_ __dut__._2325_/A __dut__._2315_/B VGND VGND VPWR VPWR __dut__._2315_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2246_ __dut__._2246_/A1 __dut__._2246_/A2 __dut__._2245_/X VGND VGND VPWR
+ VPWR __dut__._2246_/X sky130_fd_sc_hd__a21o_4
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2177_ __dut__._2189_/A __dut__._2177_/B VGND VGND VPWR VPWR __dut__._2177_/X
+ sky130_fd_sc_hd__and2_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2573__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__.__uuf__._2274__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_138_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1917__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1549__A __dut__.__uuf__._1549_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1890__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2748__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_227_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1642__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2483__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1501_ __dut__.__uuf__._1501_/A VGND VGND VPWR VPWR __dut__.__uuf__._1501_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_117_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1432_ __dut__.__uuf__._1431_/Y __dut__.__uuf__._1423_/X __dut__.__uuf__._1322_/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._1432_/X sky130_fd_sc_hd__o21a_4
XANTENNA_clkbuf_2_2_0_tck_A clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1827__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1363_ __dut__.__uuf__._1378_/A VGND VGND VPWR VPWR __dut__.__uuf__._1363_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._3017__CLK clkbuf_5_6_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1294_ __dut__.__uuf__._1294_/A VGND VGND VPWR VPWR __dut__.__uuf__._1294_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_112_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2658__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._3080_ __dut__._3093_/CLK __dut__._3080_/D __dut__._2538_/Y VGND VGND VPWR
+ VPWR __dut__._3080_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2100_ __dut__._2100_/A1 prod[32] __dut__._2099_/X VGND VGND VPWR VPWR __dut__._3107_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2031_ __dut__._2207_/A __dut__._3072_/Q VGND VGND VPWR VPWR __dut__._2031_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2297__CLK __dut__.__uuf__._2303_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2393__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2933_ clkbuf_5_9_0_tck/X __dut__._2933_/D __dut__._2685_/Y VGND VGND VPWR
+ VPWR __dut__._2933_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2864_ __dut__._2961_/CLK __dut__._2864_/D __dut__._2754_/Y VGND VGND VPWR
+ VPWR __dut__._2864_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1737__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1815_ __dut__._1817_/A __dut__._2964_/Q VGND VGND VPWR VPWR __dut__._1815_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2795_ rst VGND VGND VPWR VPWR __dut__._2795_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1746_ __dut__._1942_/A1 tie[25] __dut__._1745_/X VGND VGND VPWR VPWR __dut__._2930_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_4_0_tck_A clkbuf_4_5_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1677_ __dut__._1891_/A __dut__._2895_/Q VGND VGND VPWR VPWR __dut__._1677_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2568__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_1_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1624__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2229_ __dut__._2325_/A __dut__._2229_/B VGND VGND VPWR VPWR __dut__._2229_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_146_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1647__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_177_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2104__A2 prod[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1981_ __dut__._2235_/B __dut__._2117_/B __dut__.__uuf__._1980_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1982_/C sky130_fd_sc_hd__o21ai_4
XFILLER_51_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1742__A __dut__.__uuf__._1904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1415_ __dut__.__uuf__._1403_/X __dut__.__uuf__._1413_/X __dut__._2309_/B
+ __dut__.__uuf__._1414_/X VGND VGND VPWR VPWR __dut__._2308_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1346_ __dut__._2337_/B VGND VGND VPWR VPWR __dut__.__uuf__._1346_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1600_ __dut__._1374_/Y mp[28] __dut__._1599_/X VGND VGND VPWR VPWR __dut__._1600_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._1189__A __dut__.__uuf__._1480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2580_ rst VGND VGND VPWR VPWR __dut__._2580_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1531_ __dut__._2509_/A __dut__._2849_/Q VGND VGND VPWR VPWR __dut__._1531_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1277_ __dut__._2363_/B VGND VGND VPWR VPWR __dut__.__uuf__._1277_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1462_ __dut__._1474_/A1 __dut__._1460_/X __dut__._1461_/X VGND VGND VPWR
+ VPWR __dut__._2831_/D sky130_fd_sc_hd__a21o_4
XFILLER_37_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1393_ __dut__._2189_/A __dut__._2813_/Q VGND VGND VPWR VPWR __dut__._1393_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3063_ clkbuf_5_6_0_tck/X __dut__._3063_/D __dut__._2555_/Y VGND VGND VPWR
+ VPWR __dut__._3063_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2014_ __dut__._2014_/A1 tie[159] __dut__._2013_/X VGND VGND VPWR VPWR __dut__._3064_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_41_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpsn_inst_psn_buff_0 __dut__._1373_/Y VGND VGND VPWR VPWR psn_inst_psn_buff_9/A sky130_fd_sc_hd__buf_8
XFILLER_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_272_ _290_/CLK _272_/D VGND VGND VPWR VPWR _272_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_psn_inst_psn_buff_30_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2916_ clkbuf_5_9_0_tck/X __dut__._2916_/D __dut__._2702_/Y VGND VGND VPWR
+ VPWR __dut__._2916_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2847_ __dut__._2941_/CLK __dut__._2847_/D __dut__._2771_/Y VGND VGND VPWR
+ VPWR __dut__._2847_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1467__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2778_ rst VGND VGND VPWR VPWR __dut__._2778_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_1_0___dut__.__uuf__.__clk_source___A clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1729_ __dut__._2189_/A __dut__._2921_/Q VGND VGND VPWR VPWR __dut__._1729_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2761__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_294_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1377__A tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2180_ __dut__.__uuf__._2216_/CLK __dut__._2140_/X __dut__.__uuf__._1626_/X
+ VGND VGND VPWR VPWR __dut__._2141_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1200_ __dut__.__uuf__._1200_/A VGND VGND VPWR VPWR __dut__.__uuf__._1200_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1131_ __dut__.__uuf__._1131_/A VGND VGND VPWR VPWR __dut__.__uuf__._1131_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_102_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__273__CLK _274_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1062_ __dut__.__uuf__._1071_/A VGND VGND VPWR VPWR __dut__.__uuf__._1062_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_83_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2001__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1964_ __dut__.__uuf__._1921_/X __dut__.__uuf__._1962_/B __dut__.__uuf__._1962_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1965_/C sky130_fd_sc_hd__o21a_4
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1895_ __dut__._2203_/B __dut__._2209_/B VGND VGND VPWR VPWR __dut__.__uuf__._1896_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_149_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2671__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_40 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2126_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_152_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2701_ rst VGND VGND VPWR VPWR __dut__._2701_/Y sky130_fd_sc_hd__inv_2
Xpsn_inst_psn_buff_73 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1426_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_62 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2238_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_51 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2288_/A1
+ sky130_fd_sc_hd__buf_4
XFILLER_144_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_84 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1518_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_95 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2290_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2632_ rst VGND VGND VPWR VPWR __dut__._2632_/Y sky130_fd_sc_hd__inv_2
X__dut__._2563_ rst VGND VGND VPWR VPWR __dut__._2563_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1329_ __dut__.__uuf__._1328_/Y __dut__.__uuf__._1321_/X __dut__.__uuf__._1322_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1329_/X sky130_fd_sc_hd__o21a_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1514_ __dut__._1514_/A1 __dut__._1512_/X __dut__._1513_/X VGND VGND VPWR
+ VPWR __dut__._2844_/D sky130_fd_sc_hd__a21o_4
XFILLER_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_78_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2494_ __dut__._2502_/A1 __dut__._2494_/A2 __dut__._2493_/X VGND VGND VPWR
+ VPWR __dut__._2494_/X sky130_fd_sc_hd__a21o_4
XFILLER_64_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1445_ __dut__._1445_/A __dut__._2826_/Q VGND VGND VPWR VPWR __dut__._1445_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_74_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1376_ mc[0] __dut__._1374_/Y __dut__._1375_/X VGND VGND VPWR VPWR __dut__._1376_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_70_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3046_ __dut__._3058_/CLK __dut__._3046_/D __dut__._2572_/Y VGND VGND VPWR
+ VPWR __dut__._3046_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2004__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_255_ _306_/CLK tms VGND VGND VPWR VPWR _256_/D sky130_fd_sc_hd__dfxtp_4
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2581__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_186_ _267_/Q _187_/B VGND VGND VPWR VPWR _266_/D sky130_fd_sc_hd__or2_4
XFILLER_142_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1925__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_1_0_tck_A clkbuf_3_1_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2756__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2208__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1680_ __dut__.__uuf__._1680_/A __dut__.__uuf__._1680_/B __dut__.__uuf__._1680_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1681_/A sky130_fd_sc_hd__or3_4
XFILLER_146_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2491__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2301_ __dut__.__uuf__._2303_/CLK __dut__._2382_/X __dut__.__uuf__._1213_/X
+ VGND VGND VPWR VPWR prod[0] sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_4_12_0_tck_A clkbuf_3_6_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2232_ __dut__.__uuf__._2240_/CLK __dut__._2244_/X __dut__.__uuf__._1553_/X
+ VGND VGND VPWR VPWR __dut__._2245_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_141_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1835__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2163_ __dut__.__uuf__._2303_/CLK __dut__._2106_/X __dut__.__uuf__._1646_/X
+ VGND VGND VPWR VPWR __dut__._2107_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_87_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2094_ VGND VGND VPWR VPWR __dut__.__uuf__._2094_/HI tie[101] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1114_ __dut__.__uuf__._1464_/A VGND VGND VPWR VPWR __dut__.__uuf__._1173_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_68_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1045_ __dut__.__uuf__._1992_/A VGND VGND VPWR VPWR __dut__.__uuf__._1056_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2482__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2666__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1947_ __dut__.__uuf__._1940_/A __dut__.__uuf__._1945_/B __dut__.__uuf__._1936_/X
+ VGND VGND VPWR VPWR __dut__._2218_/A2 sky130_fd_sc_hd__o21a_4
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1878_ __dut__.__uuf__._1878_/A VGND VGND VPWR VPWR __dut__.__uuf__._1880_/B
+ sky130_fd_sc_hd__inv_2
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1994_ __dut__._2004_/A1 tie[149] __dut__._1993_/X VGND VGND VPWR VPWR __dut__._3054_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_124_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2895__CLK __dut__._3106_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2615_ rst VGND VGND VPWR VPWR __dut__._2615_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1745__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2546_ rst VGND VGND VPWR VPWR __dut__._2546_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2477_ __dut__._2491_/A prod[47] VGND VGND VPWR VPWR __dut__._2477_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2576__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1428_ __dut__._1374_/Y mc[21] __dut__._1427_/X VGND VGND VPWR VPWR __dut__._1428_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_307_ _315_/CLK _307_/D trst VGND VGND VPWR VPWR _307_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._3029_ clkbuf_5_1_0_tck/X __dut__._3029_/D __dut__._2589_/Y VGND VGND VPWR
+ VPWR __dut__._3029_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_238_ _238_/A _238_/B _300_/Q _238_/D VGND VGND VPWR VPWR _239_/C sky130_fd_sc_hd__and4_4
XFILLER_11_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_169_ _281_/Q _173_/B VGND VGND VPWR VPWR _280_/D sky130_fd_sc_hd__and2_4
XFILLER_112_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1655__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3050__CLK __dut__._3058_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_257_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2464__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2180__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_53_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1801_ __dut__.__uuf__._1844_/A __dut__.__uuf__._1801_/B __dut__.__uuf__._1801_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1802_/A sky130_fd_sc_hd__or3_4
XFILLER_21_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1732_ __dut__._1624_/X VGND VGND VPWR VPWR __dut__.__uuf__._1736_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_147_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1663_ __dut__._2367_/B __dut__._1472_/X VGND VGND VPWR VPWR __dut__.__uuf__._1663_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_146_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1594_ __dut__.__uuf__._1596_/A VGND VGND VPWR VPWR __dut__.__uuf__._1594_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_102_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2215_ __dut__.__uuf__._2225_/CLK __dut__._2210_/X __dut__.__uuf__._1583_/X
+ VGND VGND VPWR VPWR __dut__._2211_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2400_ __dut__._2412_/A1 __dut__._2400_/A2 __dut__._2399_/X VGND VGND VPWR
+ VPWR __dut__._2400_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2146_ VGND VGND VPWR VPWR __dut__.__uuf__._2146_/HI tie[153] sky130_fd_sc_hd__conb_1
XFILLER_69_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2331_ __dut__._2407_/A __dut__._2331_/B VGND VGND VPWR VPWR __dut__._2331_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._2077_ VGND VGND VPWR VPWR __dut__.__uuf__._2077_/HI tie[84] sky130_fd_sc_hd__conb_1
XFILLER_84_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2262_ __dut__._2262_/A1 __dut__._2262_/A2 __dut__._2261_/X VGND VGND VPWR
+ VPWR __dut__._2262_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1028_ __dut__.__uuf__._1074_/A VGND VGND VPWR VPWR __dut__.__uuf__._1603_/A
+ sky130_fd_sc_hd__buf_2
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2193_ __dut__._2197_/A __dut__._2193_/B VGND VGND VPWR VPWR __dut__._2193_/X
+ sky130_fd_sc_hd__and2_4
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_205 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2005_/A sky130_fd_sc_hd__buf_4
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_227 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2417_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_216 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2095_/A sky130_fd_sc_hd__buf_2
XFILLER_129_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpsn_inst_psn_buff_249 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1589_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_238 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1801_/A sky130_fd_sc_hd__buf_2
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1977_ __dut__._2005_/A __dut__._3045_/Q VGND VGND VPWR VPWR __dut__._1977_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_4_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._3073__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1475__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2529_ rst VGND VGND VPWR VPWR __dut__._2529_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1385__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2000_ VGND VGND VPWR VPWR __dut__.__uuf__._2000_/HI tie[7] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._1488__A2 mp[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1715_ __dut__.__uuf__._1736_/A __dut__.__uuf__._1715_/B __dut__.__uuf__._1715_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1716_/A sky130_fd_sc_hd__or3_4
XANTENNA___dut__._1412__A2 mc[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1480__A __dut__.__uuf__._1480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1900_ __dut__._2004_/A1 tie[102] __dut__._1899_/X VGND VGND VPWR VPWR __dut__._3007_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2880_ __dut__._3106_/CLK __dut__._2880_/D __dut__._2738_/Y VGND VGND VPWR
+ VPWR __dut__._2880_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1646_ __dut__.__uuf__._1992_/A VGND VGND VPWR VPWR __dut__.__uuf__._1646_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1577_ __dut__.__uuf__._1578_/A VGND VGND VPWR VPWR __dut__.__uuf__._1577_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1831_ __dut__._2507_/A __dut__._2972_/Q VGND VGND VPWR VPWR __dut__._1831_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_150_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1762_ __dut__._1780_/A1 tie[33] __dut__._1761_/X VGND VGND VPWR VPWR __dut__._2938_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1693_ __dut__._1817_/A __dut__._2903_/Q VGND VGND VPWR VPWR __dut__._1693_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2933__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2129_ VGND VGND VPWR VPWR __dut__.__uuf__._2129_/HI tie[136] sky130_fd_sc_hd__conb_1
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2314_ __dut__._2318_/A1 __dut__._2314_/A2 __dut__._2313_/X VGND VGND VPWR
+ VPWR __dut__._2314_/X sky130_fd_sc_hd__a21o_4
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_60_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2245_ __dut__._2245_/A __dut__._2245_/B VGND VGND VPWR VPWR __dut__._2245_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2176_ __dut__._2184_/A1 __dut__._2176_/A2 __dut__._2175_/X VGND VGND VPWR
+ VPWR __dut__._2176_/X sky130_fd_sc_hd__a21o_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1933__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_122_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2764__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1500_ __dut__.__uuf__._1486_/X __dut__.__uuf__._1480_/X __dut__._2271_/B
+ __dut__.__uuf__._1491_/X __dut__.__uuf__._1499_/X VGND VGND VPWR VPWR __dut__._2270_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_144_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1431_ __dut__._2303_/B VGND VGND VPWR VPWR __dut__.__uuf__._1431_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_132_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1362_ __dut__.__uuf__._1361_/Y __dut__.__uuf__._1347_/X __dut__.__uuf__._1348_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1362_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1293_ __dut__.__uuf__._1709_/A VGND VGND VPWR VPWR __dut__.__uuf__._1294_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_131_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2030_ __dut__._2030_/A1 tie[167] __dut__._2029_/X VGND VGND VPWR VPWR __dut__._3072_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_81_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2674__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2932_ clkbuf_5_0_0_tck/X __dut__._2932_/D __dut__._2686_/Y VGND VGND VPWR
+ VPWR __dut__._2932_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1629_ __dut__.__uuf__._1633_/A VGND VGND VPWR VPWR __dut__.__uuf__._1629_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2863_ __dut__._2961_/CLK __dut__._2863_/D __dut__._2755_/Y VGND VGND VPWR
+ VPWR __dut__._2863_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1814_ __dut__._1816_/A1 tie[59] __dut__._1813_/X VGND VGND VPWR VPWR __dut__._2964_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2794_ rst VGND VGND VPWR VPWR __dut__._2794_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1745_ __dut__._2189_/A __dut__._2929_/Q VGND VGND VPWR VPWR __dut__._1745_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_89_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1753__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1676_ __dut__._2502_/A1 prod[55] __dut__._1675_/X VGND VGND VPWR VPWR __dut__._2895_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_67_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1624__A2 mc[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2228_ __dut__._2228_/A1 __dut__._2228_/A2 __dut__._2227_/X VGND VGND VPWR
+ VPWR __dut__._2228_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2584__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2159_ __dut__._2207_/A __dut__._2159_/B VGND VGND VPWR VPWR __dut__._2159_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1388__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1560__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1663__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2759__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1980_ __dut__.__uuf__._1980_/A VGND VGND VPWR VPWR __dut__.__uuf__._1980_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_63_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1414_ __dut__.__uuf__._1414_/A VGND VGND VPWR VPWR __dut__.__uuf__._1414_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1345_ __dut__.__uuf__._1360_/A VGND VGND VPWR VPWR __dut__.__uuf__._1345_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1530_ __dut__._1562_/A1 __dut__._1528_/X __dut__._1529_/X VGND VGND VPWR
+ VPWR __dut__._2848_/D sky130_fd_sc_hd__a21o_4
XFILLER_113_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2669__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1276_ __dut__.__uuf__._1280_/A VGND VGND VPWR VPWR __dut__.__uuf__._1276_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1461_ __dut__._2325_/A __dut__._2830_/Q VGND VGND VPWR VPWR __dut__._1461_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1392_ __dut__._1374_/Y mc[13] __dut__._1391_/X VGND VGND VPWR VPWR __dut__._1392_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2264__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._3062_ clkbuf_5_6_0_tck/X __dut__._3062_/D __dut__._2556_/Y VGND VGND VPWR
+ VPWR __dut__._3062_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2013_ __dut__._2207_/A __dut__._3063_/Q VGND VGND VPWR VPWR __dut__._2013_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_1 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1932_/A1 sky130_fd_sc_hd__buf_2
X_271_ _271_/CLK _271_/D VGND VGND VPWR VPWR _271_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_23_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2915_ clkbuf_5_9_0_tck/X __dut__._2915_/D __dut__._2703_/Y VGND VGND VPWR
+ VPWR __dut__._2915_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2846_ __dut__._2846_/CLK __dut__._2846_/D __dut__._2772_/Y VGND VGND VPWR
+ VPWR __dut__._2846_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2777_ rst VGND VGND VPWR VPWR __dut__._2777_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1728_ __dut__._1760_/A1 tie[16] __dut__._1727_/X VGND VGND VPWR VPWR __dut__._2921_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1483__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2098__A2 prod[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2579__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1659_ __dut__._2491_/A __dut__._2886_/Q VGND VGND VPWR VPWR __dut__._1659_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_94_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3007__CLK _274_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_287_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1377__B __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1130_ __dut__.__uuf__._1118_/X __dut__.__uuf__._1129_/X prod[29]
+ prod[30] __dut__.__uuf__._1126_/X VGND VGND VPWR VPWR __dut__._2440_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1393__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2489__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1061_ __dut__.__uuf__._1057_/X __dut__.__uuf__._1054_/X prod[52]
+ prod[53] __dut__.__uuf__._1051_/X VGND VGND VPWR VPWR __dut__._2486_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_56_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1963_ __dut__.__uuf__._1963_/A VGND VGND VPWR VPWR __dut__.__uuf__._1965_/B
+ sky130_fd_sc_hd__inv_2
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1894_ __dut__._1432_/X VGND VGND VPWR VPWR __dut__.__uuf__._1898_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_30 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2148_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_152_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_41 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2332_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_74 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1414_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2700_ rst VGND VGND VPWR VPWR __dut__._2700_/Y sky130_fd_sc_hd__inv_2
Xpsn_inst_psn_buff_63 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2246_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_52 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2310_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1524__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_85 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1522_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2631_ rst VGND VGND VPWR VPWR __dut__._2631_/Y sky130_fd_sc_hd__inv_2
Xpsn_inst_psn_buff_96 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2296_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2562_ rst VGND VGND VPWR VPWR __dut__._2562_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2399__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1328_ __dut__._2345_/B VGND VGND VPWR VPWR __dut__.__uuf__._1328_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1513_ __dut__._2189_/A __dut__._2842_/Q VGND VGND VPWR VPWR __dut__._1513_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2493_ __dut__._2497_/A prod[55] VGND VGND VPWR VPWR __dut__._2493_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1647__B __dut__._2109_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1259_ __dut__._2367_/B VGND VGND VPWR VPWR __dut__.__uuf__._1703_/A
+ sky130_fd_sc_hd__inv_2
X__dut__._1444_ __dut__._1374_/Y mc[25] __dut__._1443_/X VGND VGND VPWR VPWR __dut__._1444_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_86_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1375_ __dut__._2810_/Q __dut__._2509_/A VGND VGND VPWR VPWR __dut__._1375_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_82_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3045_ __dut__._3058_/CLK __dut__._3045_/D __dut__._2573_/Y VGND VGND VPWR
+ VPWR __dut__._3045_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_254_ _199_/A _307_/Q VGND VGND VPWR VPWR _254_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_185_ _268_/Q _187_/B VGND VGND VPWR VPWR _267_/D sky130_fd_sc_hd__or2_4
XFILLER_142_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2829_ __dut__._2836_/CLK __dut__._2829_/D __dut__._2789_/Y VGND VGND VPWR
+ VPWR __dut__._2829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1941__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_202_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2772__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2300_ __dut__.__uuf__._2303_/CLK __dut__._2380_/X __dut__.__uuf__._1216_/X
+ VGND VGND VPWR VPWR __dut__._2381_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2231_ __dut__.__uuf__._2240_/CLK __dut__._2242_/X __dut__.__uuf__._1556_/X
+ VGND VGND VPWR VPWR __dut__._2243_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2162_ VGND VGND VPWR VPWR __dut__.__uuf__._2162_/HI tie[169] sky130_fd_sc_hd__conb_1
XFILLER_125_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2093_ VGND VGND VPWR VPWR __dut__.__uuf__._2093_/HI tie[100] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1113_ __dut__.__uuf__._1117_/A VGND VGND VPWR VPWR __dut__.__uuf__._1113_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1044_ __dut__.__uuf__._1043_/X __dut__.__uuf__._1040_/X prod[58]
+ prod[59] __dut__.__uuf__._1036_/X VGND VGND VPWR VPWR __dut__._2498_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._2302__CLK __dut__.__uuf__._2303_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1946_ __dut__.__uuf__._1946_/A VGND VGND VPWR VPWR __dut__._2220_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2682__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1877_ __dut__.__uuf__._1898_/A __dut__.__uuf__._1877_/B __dut__.__uuf__._1877_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1878_/A sky130_fd_sc_hd__or3_4
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1993_ __dut__._2005_/A __dut__._3053_/Q VGND VGND VPWR VPWR __dut__._1993_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_137_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2614_ rst VGND VGND VPWR VPWR __dut__._2614_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2170__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2545_ rst VGND VGND VPWR VPWR __dut__._2545_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_90_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1761__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2476_ __dut__._2488_/A1 __dut__._2476_/A2 __dut__._2475_/X VGND VGND VPWR
+ VPWR __dut__._2476_/X sky130_fd_sc_hd__a21o_4
XFILLER_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1427_ __dut__._2509_/A __dut__._2823_/Q VGND VGND VPWR VPWR __dut__._1427_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_131_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1984__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2592__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._3028_ clkbuf_5_1_0_tck/X __dut__._3028_/D __dut__._2590_/Y VGND VGND VPWR
+ VPWR __dut__._3028_/Q sky130_fd_sc_hd__dfrtp_4
X_306_ _306_/CLK _306_/D trst VGND VGND VPWR VPWR _306_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_42_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_237_ _237_/A _313_/Q VGND VGND VPWR VPWR _238_/D sky130_fd_sc_hd__nor2_4
XFILLER_143_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_168_ _282_/Q _173_/B VGND VGND VPWR VPWR _281_/D sky130_fd_sc_hd__and2_4
XFILLER_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2767__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_152_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1671__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1800_ __dut__._2167_/B __dut__._2173_/B __dut__.__uuf__._1799_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1801_/C sky130_fd_sc_hd__o21ai_4
XFILLER_34_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1731_ __dut__.__uuf__._1724_/A __dut__.__uuf__._1729_/B __dut__.__uuf__._1720_/X
+ VGND VGND VPWR VPWR __dut__._2138_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_21_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1662_ __dut__.__uuf__._1654_/A __dut__.__uuf__._1659_/B __dut__.__uuf__._1661_/X
+ VGND VGND VPWR VPWR __dut__._2110_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_119_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2007__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1593_ __dut__.__uuf__._1596_/A VGND VGND VPWR VPWR __dut__.__uuf__._1593_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_106_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2214_ __dut__.__uuf__._2216_/CLK __dut__._2208_/X __dut__.__uuf__._1584_/X
+ VGND VGND VPWR VPWR __dut__._2209_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2145_ VGND VGND VPWR VPWR __dut__.__uuf__._2145_/HI tie[152] sky130_fd_sc_hd__conb_1
XFILLER_130_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2330_ __dut__._2332_/A1 __dut__._2330_/A2 __dut__._2329_/X VGND VGND VPWR
+ VPWR __dut__._2330_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2677__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2076_ VGND VGND VPWR VPWR __dut__.__uuf__._2076_/HI tie[83] sky130_fd_sc_hd__conb_1
XFILLER_44_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2261_ __dut__._2261_/A __dut__._2261_/B VGND VGND VPWR VPWR __dut__._2261_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1027_ rst VGND VGND VPWR VPWR __dut__.__uuf__._1074_/A sky130_fd_sc_hd__inv_2
XFILLER_43_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2192_ __dut__._2192_/A1 __dut__._2192_/A2 __dut__._2191_/X VGND VGND VPWR
+ VPWR __dut__._2192_/X sky130_fd_sc_hd__a21o_4
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__286__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_206 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1969_/A sky130_fd_sc_hd__buf_2
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_217 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2435_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_228 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2069_/A sky130_fd_sc_hd__buf_2
XFILLER_101_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1966__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_239 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1803_/A sky130_fd_sc_hd__buf_2
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1929_ __dut__.__uuf__._1929_/A VGND VGND VPWR VPWR __dut__.__uuf__._1929_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1976_ __dut__._2004_/A1 tie[140] __dut__._1975_/X VGND VGND VPWR VPWR __dut__._3045_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_125_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2528_ rst VGND VGND VPWR VPWR __dut__._2528_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2587__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__299__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1491__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2459_ __dut__._2491_/A prod[38] VGND VGND VPWR VPWR __dut__._2459_/X sky130_fd_sc_hd__and2_4
XFILLER_62_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2382__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2885__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1948__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1714_ __dut__._2135_/B __dut__._2141_/B __dut__.__uuf__._1713_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1715_/C sky130_fd_sc_hd__o21ai_4
XFILLER_119_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1645_ __dut__.__uuf__._1645_/A VGND VGND VPWR VPWR __dut__.__uuf__._1645_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_107_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1830_ __dut__._1830_/A1 tie[67] __dut__._1829_/X VGND VGND VPWR VPWR __dut__._2972_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1576_ __dut__.__uuf__._1578_/A VGND VGND VPWR VPWR __dut__.__uuf__._1576_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1761_ __dut__._2189_/A __dut__._2937_/Q VGND VGND VPWR VPWR __dut__._1761_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1692_ __dut__._2412_/A1 prod[63] __dut__._1691_/X VGND VGND VPWR VPWR __dut__._2903_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2128_ VGND VGND VPWR VPWR __dut__.__uuf__._2128_/HI tie[135] sky130_fd_sc_hd__conb_1
XANTENNA___dut__.__uuf__._1936__A __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2059_ VGND VGND VPWR VPWR __dut__.__uuf__._2059_/HI tie[66] sky130_fd_sc_hd__conb_1
X__dut__._2313_ __dut__._2325_/A __dut__._2313_/B VGND VGND VPWR VPWR __dut__._2313_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2244_ __dut__._2246_/A1 __dut__._2244_/A2 __dut__._2243_/X VGND VGND VPWR
+ VPWR __dut__._2244_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2175_ __dut__._2189_/A __dut__._2175_/B VGND VGND VPWR VPWR __dut__._2175_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2364__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1959_ __dut__._2207_/A __dut__._3036_/Q VGND VGND VPWR VPWR __dut__._1959_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2170__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_97_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1933__B __dut__._3023_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_115_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2780__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1430_ __dut__.__uuf__._1434_/A VGND VGND VPWR VPWR __dut__.__uuf__._1430_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_144_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1361_ __dut__._2331_/B VGND VGND VPWR VPWR __dut__.__uuf__._1361_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_132_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1292_ __dut__.__uuf__._1292_/A VGND VGND VPWR VPWR __dut__.__uuf__._1709_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_86_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_tck clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR clkbuf_3_7_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_66_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._3063__CLK clkbuf_5_6_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1491__A __dut__.__uuf__._1533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2931_ clkbuf_5_0_0_tck/X __dut__._2931_/D __dut__._2687_/Y VGND VGND VPWR
+ VPWR __dut__._2931_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2690__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2193__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1628_ __dut__.__uuf__._1628_/A VGND VGND VPWR VPWR __dut__.__uuf__._1633_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2346__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2862_ __dut__._2961_/CLK __dut__._2862_/D __dut__._2756_/Y VGND VGND VPWR
+ VPWR __dut__._2862_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1813_ __dut__._1817_/A __dut__._2963_/Q VGND VGND VPWR VPWR __dut__._1813_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2793_ rst VGND VGND VPWR VPWR __dut__._2793_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1559_ __dut__.__uuf__._1562_/A VGND VGND VPWR VPWR __dut__.__uuf__._1559_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_122_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1744_ __dut__._1942_/A1 tie[24] __dut__._1743_/X VGND VGND VPWR VPWR __dut__._2929_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_150_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1675_ __dut__._2491_/A __dut__._2894_/Q VGND VGND VPWR VPWR __dut__._1675_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_83_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2227_ __dut__._2325_/A __dut__._2227_/B VGND VGND VPWR VPWR __dut__._2227_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_83_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_5_0___dut__.__uuf__.__clk_source__ clkbuf_4_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2225_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__._2158_ __dut__._2172_/A1 __dut__._2158_/A2 __dut__._2157_/X VGND VGND VPWR
+ VPWR __dut__._2158_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1388__A2 mc[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2089_ __dut__._2431_/A __dut__._3101_/Q VGND VGND VPWR VPWR __dut__._2089_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_9_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1560__A2 mp[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3086__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_232_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2775__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2923__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2328__A1 __dut__._2332_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1413_ __dut__.__uuf__._1412_/Y __dut__.__uuf__._1398_/X __dut__.__uuf__._1399_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1413_/X sky130_fd_sc_hd__o21a_4
XFILLER_144_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2015__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1344_ __dut__.__uuf__._1338_/X __dut__.__uuf__._1343_/X __dut__._2337_/B
+ __dut__.__uuf__._1338_/X VGND VGND VPWR VPWR __dut__._2336_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1275_ __dut__.__uuf__._1271_/X __dut__.__uuf__._1274_/X __dut__._2363_/B
+ __dut__.__uuf__._1271_/X VGND VGND VPWR VPWR __dut__._2362_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1486__A __dut__.__uuf__._1549_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2500__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1460_ __dut__._1374_/Y mc[29] __dut__._1459_/X VGND VGND VPWR VPWR __dut__._1460_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_58_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1391_ __dut__._2509_/A __dut__._2814_/Q VGND VGND VPWR VPWR __dut__._1391_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_37_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2685__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._3061_ clkbuf_5_6_0_tck/X __dut__._3061_/D __dut__._2557_/Y VGND VGND VPWR
+ VPWR __dut__._3061_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2012_ __dut__._2012_/A1 tie[158] __dut__._2011_/X VGND VGND VPWR VPWR __dut__._3063_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpsn_inst_psn_buff_2 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1930_/A1 sky130_fd_sc_hd__buf_2
XFILLER_139_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_270_ _271_/CLK _270_/D VGND VGND VPWR VPWR _270_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__255__D tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_16_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2914_ clkbuf_5_9_0_tck/X __dut__._2914_/D __dut__._2704_/Y VGND VGND VPWR
+ VPWR __dut__._2914_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2845_ __dut__._2846_/CLK __dut__._2845_/D __dut__._2773_/Y VGND VGND VPWR
+ VPWR __dut__._2845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2776_ rst VGND VGND VPWR VPWR __dut__._2776_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1727_ __dut__._2189_/A __dut__._2920_/Q VGND VGND VPWR VPWR __dut__._1727_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1658_ __dut__._2488_/A1 prod[46] __dut__._1657_/X VGND VGND VPWR VPWR __dut__._2886_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1589_ __dut__._1589_/A __dut__._2862_/Q VGND VGND VPWR VPWR __dut__._1589_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2595__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1939__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1196__A3 prod[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1060_ __dut__.__uuf__._1071_/A VGND VGND VPWR VPWR __dut__.__uuf__._1060_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1962_ __dut__.__uuf__._1982_/A __dut__.__uuf__._1962_/B __dut__.__uuf__._1962_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1963_/A sky130_fd_sc_hd__or3_4
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1893_ __dut__.__uuf__._1886_/A __dut__.__uuf__._1891_/B __dut__.__uuf__._1882_/X
+ VGND VGND VPWR VPWR __dut__._2198_/A2 sky130_fd_sc_hd__o21a_4
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3101__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_20 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2014_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_31 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2142_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_42 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2228_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_64 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1446_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_53 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2308_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_75 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1390_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2630_ rst VGND VGND VPWR VPWR __dut__._2630_/Y sky130_fd_sc_hd__inv_2
Xpsn_inst_psn_buff_86 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1526_/A1 sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1524__A2 mp[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_97 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2300_/A1 sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1327_ __dut__.__uuf__._1378_/A VGND VGND VPWR VPWR __dut__.__uuf__._1327_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2231__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2561_ rst VGND VGND VPWR VPWR __dut__._2561_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2399__B prod[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1512_ __dut__._1374_/Y mp[8] __dut__._1511_/X VGND VGND VPWR VPWR __dut__._1512_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._2492_ __dut__._2502_/A1 __dut__._2492_/A2 __dut__._2491_/X VGND VGND VPWR
+ VPWR __dut__._2492_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1258_ __dut__.__uuf__._1280_/A VGND VGND VPWR VPWR __dut__.__uuf__._1258_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1189_ __dut__.__uuf__._1480_/A VGND VGND VPWR VPWR __dut__.__uuf__._1189_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1443_ __dut__._2509_/A __dut__._2827_/Q VGND VGND VPWR VPWR __dut__._1443_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1374_ __dut__._2509_/A VGND VGND VPWR VPWR __dut__._1374_/Y sky130_fd_sc_hd__inv_8
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3044_ __dut__._3058_/CLK __dut__._3044_/D __dut__._2574_/Y VGND VGND VPWR
+ VPWR __dut__._3044_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1460__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_253_ _196_/X _259_/Q VGND VGND VPWR VPWR _253_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1759__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_184_ _269_/Q _191_/B VGND VGND VPWR VPWR _268_/D sky130_fd_sc_hd__and2_4
XFILLER_127_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2828_ clkbuf_5_3_0_tck/X __dut__._2828_/D __dut__._2790_/Y VGND VGND VPWR
+ VPWR __dut__._2828_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2759_ rst VGND VGND VPWR VPWR __dut__._2759_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1669__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2230_ __dut__.__uuf__._2230_/CLK __dut__._2240_/X __dut__.__uuf__._1559_/X
+ VGND VGND VPWR VPWR __dut__._2241_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2161_ VGND VGND VPWR VPWR __dut__.__uuf__._2161_/HI tie[168] sky130_fd_sc_hd__conb_1
XFILLER_130_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2092_ VGND VGND VPWR VPWR __dut__.__uuf__._2092_/HI tie[99] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1112_ __dut__.__uuf__._1103_/X __dut__.__uuf__._1099_/X prod[35]
+ prod[36] __dut__.__uuf__._1111_/X VGND VGND VPWR VPWR __dut__._2452_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1043_ __dut__.__uuf__._1088_/A VGND VGND VPWR VPWR __dut__.__uuf__._1043_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_110_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1945_ __dut__.__uuf__._1975_/A __dut__.__uuf__._1945_/B __dut__.__uuf__._1945_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1946_/A sky130_fd_sc_hd__or3_4
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1876_ __dut__._2195_/B __dut__._2201_/B __dut__.__uuf__._1875_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1877_/C sky130_fd_sc_hd__o21ai_4
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1579__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1992_ __dut__._2004_/A1 tie[148] __dut__._1991_/X VGND VGND VPWR VPWR __dut__._3053_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_109_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2613_ rst VGND VGND VPWR VPWR __dut__._2613_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2359_ __dut__.__uuf__._2364_/CLK __dut__._2498_/X __dut__.__uuf__._1042_/X
+ VGND VGND VPWR VPWR prod[58] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2203__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2544_ rst VGND VGND VPWR VPWR __dut__._2544_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_83_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2475_ __dut__._2491_/A prod[46] VGND VGND VPWR VPWR __dut__._2475_/X sky130_fd_sc_hd__and2_4
X__dut__._1426_ __dut__._1426_/A1 __dut__._1424_/X __dut__._1425_/X VGND VGND VPWR
+ VPWR __dut__._2822_/D sky130_fd_sc_hd__a21o_4
XFILLER_62_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_305_ _313_/CLK _305_/D trst VGND VGND VPWR VPWR _305_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._2277__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._3027_ clkbuf_5_1_0_tck/X __dut__._3027_/D __dut__._2591_/Y VGND VGND VPWR
+ VPWR __dut__._3027_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_236_ _305_/Q _306_/Q VGND VGND VPWR VPWR _236_/Y sky130_fd_sc_hd__nor2_4
XFILLER_156_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_167_ _283_/Q _172_/B VGND VGND VPWR VPWR _282_/D sky130_fd_sc_hd__or2_4
XFILLER_112_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2113__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1672__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_145_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1424__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2783__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1730_ __dut__.__uuf__._1730_/A VGND VGND VPWR VPWR __dut__._2140_/A2
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1399__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1661_ __dut__.__uuf__._1828_/A VGND VGND VPWR VPWR __dut__.__uuf__._1661_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1592_ __dut__.__uuf__._1596_/A VGND VGND VPWR VPWR __dut__.__uuf__._1592_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__.__uuf__._1759__A __dut__.__uuf__._1982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2023__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2213_ __dut__.__uuf__._2216_/CLK __dut__._2206_/X __dut__.__uuf__._1586_/X
+ VGND VGND VPWR VPWR __dut__._2207_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2144_ VGND VGND VPWR VPWR __dut__.__uuf__._2144_/HI tie[151] sky130_fd_sc_hd__conb_1
XFILLER_102_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_9_0_tck clkbuf_5_9_0_tck/A VGND VGND VPWR VPWR clkbuf_5_9_0_tck/X sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2075_ VGND VGND VPWR VPWR __dut__.__uuf__._2075_/HI tie[82] sky130_fd_sc_hd__conb_1
XFILLER_84_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2260_ __dut__._2262_/A1 __dut__._2260_/A2 __dut__._2259_/X VGND VGND VPWR
+ VPWR __dut__._2260_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1026_ __dut__.__uuf__._1019_/X __dut__.__uuf__._1023_/X prod[63]
+ __dut__._2113_/B __dut__.__uuf__._1025_/X VGND VGND VPWR VPWR __dut__._2508_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_71_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2191_ __dut__._2197_/A __dut__._2191_/B VGND VGND VPWR VPWR __dut__._2191_/X
+ sky130_fd_sc_hd__and2_4
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_207 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1967_/A sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2693__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_218 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2491_/A sky130_fd_sc_hd__buf_4
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_229 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2391_/A sky130_fd_sc_hd__buf_2
XFILLER_24_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1928_ __dut__._2215_/B __dut__._2221_/B VGND VGND VPWR VPWR __dut__.__uuf__._1929_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_101_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1859_ __dut__.__uuf__._1859_/A VGND VGND VPWR VPWR __dut__._2188_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_138_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1975_ __dut__._2005_/A __dut__._3044_/Q VGND VGND VPWR VPWR __dut__._1975_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2527_ rst VGND VGND VPWR VPWR __dut__._2527_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1654__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2458_ __dut__._2502_/A1 __dut__._2458_/A2 __dut__._2457_/X VGND VGND VPWR
+ VPWR __dut__._2458_/X sky130_fd_sc_hd__a21o_4
XFILLER_142_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1409_ __dut__._2189_/A __dut__._2817_/Q VGND VGND VPWR VPWR __dut__._1409_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2389_ __dut__._2389_/A prod[3] VGND VGND VPWR VPWR __dut__._2389_/X sky130_fd_sc_hd__and2_4
XFILLER_43_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1406__A1 __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_219_ _294_/Q _293_/Q _222_/A VGND VGND VPWR VPWR _293_/D sky130_fd_sc_hd__o21a_4
XFILLER_128_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1947__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_262_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2778__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2497__B prod[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1713_ __dut__.__uuf__._1713_/A VGND VGND VPWR VPWR __dut__.__uuf__._1713_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_119_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1644_ __dut__.__uuf__._1645_/A VGND VGND VPWR VPWR __dut__.__uuf__._1644_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1575_ __dut__.__uuf__._1578_/A VGND VGND VPWR VPWR __dut__.__uuf__._1575_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1760_ __dut__._1760_/A1 tie[32] __dut__._1759_/X VGND VGND VPWR VPWR __dut__._2937_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_88_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1691_ __dut__._2407_/A __dut__._2902_/Q VGND VGND VPWR VPWR __dut__._1691_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_102_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2688__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2127_ VGND VGND VPWR VPWR __dut__.__uuf__._2127_/HI tie[134] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2058_ VGND VGND VPWR VPWR __dut__.__uuf__._2058_/HI tie[65] sky130_fd_sc_hd__conb_1
X__dut__._2312_ __dut__._2312_/A1 __dut__._2312_/A2 __dut__._2311_/X VGND VGND VPWR
+ VPWR __dut__._2312_/X sky130_fd_sc_hd__a21o_4
XFILLER_56_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_tck tck VGND VGND VPWR VPWR clkbuf_0_tck/X sky130_fd_sc_hd__clkbuf_16
X__dut__._2243_ __dut__._2245_/A __dut__._2243_/B VGND VGND VPWR VPWR __dut__._2243_/X
+ sky130_fd_sc_hd__and2_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2174_ __dut__._2184_/A1 __dut__._2174_/A2 __dut__._2173_/X VGND VGND VPWR
+ VPWR __dut__._2174_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1958_ __dut__._1958_/A1 tie[131] __dut__._1957_/X VGND VGND VPWR VPWR __dut__._3036_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_140_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1889_ __dut__._2491_/A __dut__._3001_/Q VGND VGND VPWR VPWR __dut__._1889_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2598__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2052__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_108_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1360_ __dut__.__uuf__._1360_/A VGND VGND VPWR VPWR __dut__.__uuf__._1360_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1102__A __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1291_ __dut__._2357_/B VGND VGND VPWR VPWR __dut__.__uuf__._1291_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_39_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2930_ clkbuf_5_0_0_tck/X __dut__._2930_/D __dut__._2688_/Y VGND VGND VPWR
+ VPWR __dut__._2930_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1627_ __dut__.__uuf__._1627_/A VGND VGND VPWR VPWR __dut__.__uuf__._1627_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2861_ __dut__._2941_/CLK __dut__._2861_/D __dut__._2757_/Y VGND VGND VPWR
+ VPWR __dut__._2861_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1587__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1812_ __dut__._1816_/A1 tie[58] __dut__._1811_/X VGND VGND VPWR VPWR __dut__._2963_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1558_ __dut__.__uuf__._1549_/X __dut__.__uuf__._1544_/X __dut__._2243_/B
+ __dut__.__uuf__._1447_/A __dut__.__uuf__._1557_/X VGND VGND VPWR VPWR __dut__._2242_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._2792_ rst VGND VGND VPWR VPWR __dut__._2792_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1743_ __dut__._2189_/A __dut__._2928_/Q VGND VGND VPWR VPWR __dut__._1743_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1489_ __dut__.__uuf__._1486_/X __dut__.__uuf__._1480_/X __dut__._2277_/B
+ __dut__.__uuf__._1469_/X __dut__.__uuf__._1488_/X VGND VGND VPWR VPWR __dut__._2276_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_107_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1674_ __dut__._2488_/A1 prod[54] __dut__._1673_/X VGND VGND VPWR VPWR __dut__._2894_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_131_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2211__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2226_ __dut__._2226_/A1 __dut__._2226_/A2 __dut__._2225_/X VGND VGND VPWR
+ VPWR __dut__._2226_/X sky130_fd_sc_hd__a21o_4
X__dut__._2157_ __dut__._2207_/A __dut__._2157_/B VGND VGND VPWR VPWR __dut__._2157_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2088_ __dut__._2488_/A1 prod[26] __dut__._2087_/X VGND VGND VPWR VPWR __dut__._3101_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1497__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2875__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2121__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_225_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2791__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1412_ __dut__._2311_/B VGND VGND VPWR VPWR __dut__.__uuf__._1412_/Y
+ sky130_fd_sc_hd__inv_2
Xclkbuf_4_15_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2364_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_144_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1343_ __dut__.__uuf__._1342_/Y __dut__.__uuf__._1321_/X __dut__.__uuf__._1322_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1343_/X sky130_fd_sc_hd__o21a_4
XFILLER_144_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1274_ __dut__.__uuf__._1266_/Y __dut__.__uuf__._1985_/A __dut__.__uuf__._1268_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1274_/X sky130_fd_sc_hd__o21a_4
XFILLER_113_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2031__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1390_ __dut__._1390_/A1 __dut__._1388_/X __dut__._1389_/X VGND VGND VPWR
+ VPWR __dut__._2813_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._3030__CLK clkbuf_5_1_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3060_ clkbuf_5_4_0_tck/X __dut__._3060_/D __dut__._2558_/Y VGND VGND VPWR
+ VPWR __dut__._3060_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2011_ __dut__._2207_/A __dut__._3062_/Q VGND VGND VPWR VPWR __dut__._2011_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_42_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_3 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1928_/A1 sky130_fd_sc_hd__buf_2
XFILLER_155_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2913_ __dut__._2509_/B __dut__._2913_/D __dut__._2705_/Y VGND VGND VPWR
+ VPWR __dut__._2913_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2844_ __dut__._2846_/CLK __dut__._2844_/D __dut__._2774_/Y VGND VGND VPWR
+ VPWR __dut__._2844_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2775_ rst VGND VGND VPWR VPWR __dut__._2775_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1726_ __dut__._1726_/A1 tie[15] __dut__._1725_/X VGND VGND VPWR VPWR __dut__._2920_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_77_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1657_ __dut__._2491_/A __dut__._2885_/Q VGND VGND VPWR VPWR __dut__._1657_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1588_ __dut__._1374_/Y mp[26] __dut__._1587_/X VGND VGND VPWR VPWR __dut__._1588_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_91_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2209_ __dut__._2507_/A __dut__._2209_/B VGND VGND VPWR VPWR __dut__._2209_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_146_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_tck clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR clkbuf_3_5_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_142_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1955__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3053__CLK __dut__._3059_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_175_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2494__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2786__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2183__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1961_ __dut__._2227_/B __dut__._2233_/B __dut__.__uuf__._1960_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1962_/C sky130_fd_sc_hd__o21ai_4
X__dut__.__uuf__._1892_ __dut__.__uuf__._1892_/A VGND VGND VPWR VPWR __dut__._2200_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_10 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2034_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_21 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2012_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_117_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_32 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2144_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_43 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2226_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_65 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1442_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_54 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2312_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_76 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1394_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_87 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2262_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_98 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1610_/A1 sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1041__B1 prod[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1326_ __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR __dut__.__uuf__._1378_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._2560_ rst VGND VGND VPWR VPWR __dut__._2560_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1511_ __dut__._2509_/A __dut__._2844_/Q VGND VGND VPWR VPWR __dut__._1511_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2491_ __dut__._2491_/A prod[54] VGND VGND VPWR VPWR __dut__._2491_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1257_ __dut__.__uuf__._1340_/A VGND VGND VPWR VPWR __dut__.__uuf__._1280_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_104_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2696__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1188_ __dut__.__uuf__._1464_/A VGND VGND VPWR VPWR __dut__.__uuf__._1480_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1442_ __dut__._1442_/A1 __dut__._1440_/X __dut__._1441_/X VGND VGND VPWR
+ VPWR __dut__._2826_/D sky130_fd_sc_hd__a21o_4
XFILLER_100_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1373_ __dut__._2207_/A VGND VGND VPWR VPWR __dut__._1373_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3043_ __dut__._3058_/CLK __dut__._3043_/D __dut__._2575_/Y VGND VGND VPWR
+ VPWR __dut__._3043_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1460__A2 mc[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_252_ _197_/X _315_/Q VGND VGND VPWR VPWR _252_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ _183_/A VGND VGND VPWR VPWR _191_/B sky130_fd_sc_hd__buf_2
XFILLER_10_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2827_ __dut__._2836_/CLK __dut__._2827_/D __dut__._2791_/Y VGND VGND VPWR
+ VPWR __dut__._2827_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2758_ rst VGND VGND VPWR VPWR __dut__._2758_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2476__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1709_ __dut__._2189_/A __dut__._2911_/Q VGND VGND VPWR VPWR __dut__._1709_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2689_ rst VGND VGND VPWR VPWR __dut__._2689_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2400__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_292_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_1_0___dut__.__uuf__.__clk_source___A clkbuf_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2160_ VGND VGND VPWR VPWR __dut__.__uuf__._2160_/HI tie[167] sky130_fd_sc_hd__conb_1
XFILLER_130_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1111_ __dut__.__uuf__._1126_/A VGND VGND VPWR VPWR __dut__.__uuf__._1111_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2091_ VGND VGND VPWR VPWR __dut__.__uuf__._2091_/HI tie[98] sky130_fd_sc_hd__conb_1
XFILLER_96_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1042_ __dut__.__uuf__._1042_/A VGND VGND VPWR VPWR __dut__.__uuf__._1042_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_141_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1690__A2 prod[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1944_ __dut__.__uuf__._1921_/X __dut__.__uuf__._1942_/B __dut__.__uuf__._1942_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1945_/C sky130_fd_sc_hd__o21a_4
XFILLER_51_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1875_ __dut__.__uuf__._1875_/A VGND VGND VPWR VPWR __dut__.__uuf__._1875_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_137_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3099__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1991_ __dut__._2005_/A __dut__._3052_/Q VGND VGND VPWR VPWR __dut__._1991_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_126_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1595__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2612_ rst VGND VGND VPWR VPWR __dut__._2612_/Y sky130_fd_sc_hd__inv_2
XANTENNA__315__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2936__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2358_ __dut__.__uuf__._2358_/CLK __dut__._2496_/X __dut__.__uuf__._1046_/X
+ VGND VGND VPWR VPWR prod[57] sky130_fd_sc_hd__dfrtp_4
XFILLER_78_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2543_ rst VGND VGND VPWR VPWR __dut__._2543_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1309_ __dut__._2351_/B VGND VGND VPWR VPWR __dut__.__uuf__._1309_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2289_ __dut__.__uuf__._2291_/CLK __dut__._2358_/X __dut__.__uuf__._1280_/X
+ VGND VGND VPWR VPWR __dut__._2359_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2458__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_76_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2474_ __dut__._2488_/A1 __dut__._2474_/A2 __dut__._2473_/X VGND VGND VPWR
+ VPWR __dut__._2474_/X sky130_fd_sc_hd__a21o_4
XFILLER_74_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1425_ __dut__._1429_/A __dut__._2820_/Q VGND VGND VPWR VPWR __dut__._1425_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_131_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3026_ clkbuf_5_1_0_tck/X __dut__._3026_/D __dut__._2592_/Y VGND VGND VPWR
+ VPWR __dut__._3026_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_304_ _306_/CLK _304_/D trst VGND VGND VPWR VPWR _304_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_235_ _251_/Q VGND VGND VPWR VPWR tdo_paden_o sky130_fd_sc_hd__inv_2
XFILLER_156_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_166_ _284_/Q _173_/B VGND VGND VPWR VPWR _283_/D sky130_fd_sc_hd__and2_4
XFILLER_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2113__B __dut__._2113_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_138_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1424__A2 mc[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1660_ __dut__.__uuf__._1660_/A VGND VGND VPWR VPWR __dut__._2112_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_147_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1591_ __dut__.__uuf__._1597_/A VGND VGND VPWR VPWR __dut__.__uuf__._1596_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_146_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2212_ __dut__.__uuf__._2216_/CLK __dut__._2204_/X __dut__.__uuf__._1587_/X
+ VGND VGND VPWR VPWR __dut__._2205_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2143_ VGND VGND VPWR VPWR __dut__.__uuf__._2143_/HI tie[150] sky130_fd_sc_hd__conb_1
XFILLER_142_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._2074_ VGND VGND VPWR VPWR __dut__.__uuf__._2074_/HI tie[81] sky130_fd_sc_hd__conb_1
XFILLER_29_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1025_ __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR __dut__.__uuf__._1025_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2190_ __dut__._2192_/A1 __dut__._2190_/A2 __dut__._2189_/X VGND VGND VPWR
+ VPWR __dut__._2190_/X sky130_fd_sc_hd__a21o_4
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_219 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2431_/A sky130_fd_sc_hd__buf_2
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_208 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1965_/A sky130_fd_sc_hd__buf_2
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1927_ __dut__._1444_/X VGND VGND VPWR VPWR __dut__.__uuf__._1931_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_101_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1858_ __dut__.__uuf__._1869_/A __dut__.__uuf__._1858_/B __dut__.__uuf__._1858_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1859_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1789_ __dut__._2163_/B __dut__._2169_/B __dut__.__uuf__._1788_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1790_/C sky130_fd_sc_hd__o21ai_4
X__dut__._1974_ __dut__._2004_/A1 tie[139] __dut__._1973_/X VGND VGND VPWR VPWR __dut__._3044_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_125_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2526_ rst VGND VGND VPWR VPWR __dut__._2526_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2457_ __dut__._2457_/A prod[37] VGND VGND VPWR VPWR __dut__._2457_/X sky130_fd_sc_hd__and2_4
XFILLER_47_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1408_ __dut__._1374_/Y mc[17] __dut__._1407_/X VGND VGND VPWR VPWR __dut__._1408_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._2388_ __dut__._2412_/A1 __dut__._2388_/A2 __dut__._2387_/X VGND VGND VPWR
+ VPWR __dut__._2388_/X sky130_fd_sc_hd__a21o_4
XFILLER_62_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3009_ _274_/CLK __dut__._3009_/D __dut__._2609_/Y VGND VGND VPWR VPWR __dut__._3009_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_30_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_218_ _234_/A VGND VGND VPWR VPWR _222_/A sky130_fd_sc_hd__buf_2
XFILLER_144_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_149_ _239_/A _142_/Y _309_/Q _308_/Q _144_/Y VGND VGND VPWR VPWR _308_/D sky130_fd_sc_hd__a32o_4
XFILLER_143_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_255_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2794__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1712_ __dut__._2135_/B __dut__._2141_/B VGND VGND VPWR VPWR __dut__.__uuf__._1713_/A
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1643_ __dut__.__uuf__._1645_/A VGND VGND VPWR VPWR __dut__.__uuf__._1643_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1574_ __dut__.__uuf__._1578_/A VGND VGND VPWR VPWR __dut__.__uuf__._1574_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1690_ __dut__._1690_/A1 prod[62] __dut__._1689_/X VGND VGND VPWR VPWR __dut__._2902_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2126_ VGND VGND VPWR VPWR __dut__.__uuf__._2126_/HI tie[133] sky130_fd_sc_hd__conb_1
XANTENNA___dut__.__uuf__._2267__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2057_ VGND VGND VPWR VPWR __dut__.__uuf__._2057_/HI tie[64] sky130_fd_sc_hd__conb_1
XFILLER_29_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2311_ __dut__._2325_/A __dut__._2311_/B VGND VGND VPWR VPWR __dut__._2311_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2242_ __dut__._2246_/A1 __dut__._2242_/A2 __dut__._2241_/X VGND VGND VPWR
+ VPWR __dut__._2242_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1636__A2 prod[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2173_ __dut__._2189_/A __dut__._2173_/B VGND VGND VPWR VPWR __dut__._2173_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2209__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_39_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1572__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1957_ __dut__._2207_/A __dut__._3035_/Q VGND VGND VPWR VPWR __dut__._1957_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_140_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1888_ __dut__._2488_/A1 tie[96] __dut__._1887_/X VGND VGND VPWR VPWR __dut__._3001_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_97_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2509_ __dut__._2509_/A __dut__._2509_/B VGND VGND VPWR VPWR __dut__._2509_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_75_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2119__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2052__A2 prod[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_8_0_tck clkbuf_5_9_0_tck/A VGND VGND VPWR VPWR __dut__._2509_/B sky130_fd_sc_hd__clkbuf_1
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1290_ __dut__.__uuf__._1308_/A VGND VGND VPWR VPWR __dut__.__uuf__._1290_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2789__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2029__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1626_ __dut__.__uuf__._1627_/A VGND VGND VPWR VPWR __dut__.__uuf__._1626_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2860_ __dut__._2860_/CLK __dut__._2860_/D __dut__._2758_/Y VGND VGND VPWR
+ VPWR __dut__._2860_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1811_ __dut__._1817_/A __dut__._2962_/Q VGND VGND VPWR VPWR __dut__._1811_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1557_ __dut__._1484_/X __dut__.__uuf__._1550_/X __dut__._2245_/B
+ __dut__.__uuf__._1294_/A VGND VGND VPWR VPWR __dut__.__uuf__._1557_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2791_ rst VGND VGND VPWR VPWR __dut__._2791_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2699__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1742_ __dut__._1942_/A1 tie[23] __dut__._1741_/X VGND VGND VPWR VPWR __dut__._2928_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1488_ __dut__._1560_/X __dut__.__uuf__._1487_/X __dut__._2279_/B
+ __dut__.__uuf__._1470_/X VGND VGND VPWR VPWR __dut__.__uuf__._1488_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1673_ __dut__._2491_/A __dut__._2893_/Q VGND VGND VPWR VPWR __dut__._1673_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_107_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2109_ VGND VGND VPWR VPWR __dut__.__uuf__._2109_/HI tie[116] sky130_fd_sc_hd__conb_1
XFILLER_76_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2225_ __dut__._2325_/A __dut__._2225_/B VGND VGND VPWR VPWR __dut__._2225_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2156_ __dut__._2172_/A1 __dut__._2156_/A2 __dut__._2155_/X VGND VGND VPWR
+ VPWR __dut__._2156_/X sky130_fd_sc_hd__a21o_4
X__dut__._2087_ __dut__._2431_/A __dut__._3100_/Q VGND VGND VPWR VPWR __dut__._2087_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_154_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1203__A __dut__.__uuf__._1480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2989_ __dut__._3096_/CLK __dut__._2989_/D __dut__._2629_/Y VGND VGND VPWR
+ VPWR __dut__._2989_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_120_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_218_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1536__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1411_ __dut__.__uuf__._1411_/A VGND VGND VPWR VPWR __dut__.__uuf__._1411_/X
+ sky130_fd_sc_hd__buf_2
Xclkbuf_3_7_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0___dut__.__uuf__.__clk_source__/X sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1342_ __dut__._2339_/B VGND VGND VPWR VPWR __dut__.__uuf__._1342_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_104_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1273_ __dut__.__uuf__._1492_/A VGND VGND VPWR VPWR __dut__.__uuf__._1985_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2010_ __dut__._2010_/A1 tie[157] __dut__._2009_/X VGND VGND VPWR VPWR __dut__._3062_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_42_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_4 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1926_/A1 sky130_fd_sc_hd__buf_2
XFILLER_139_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2912_ __dut__._2509_/B __dut__._2912_/D __dut__._2706_/Y VGND VGND VPWR
+ VPWR __dut__._2912_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1609_ __dut__.__uuf__._1609_/A VGND VGND VPWR VPWR __dut__.__uuf__._1609_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1023__A __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2843_ clkbuf_5_3_0_tck/X __dut__._2843_/D __dut__._2775_/Y VGND VGND VPWR
+ VPWR __dut__._2843_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2774_ rst VGND VGND VPWR VPWR __dut__._2774_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1725_ __dut__._2189_/A __dut__._2919_/Q VGND VGND VPWR VPWR __dut__._1725_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1656_ __dut__._2488_/A1 prod[45] __dut__._1655_/X VGND VGND VPWR VPWR __dut__._2885_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1587_ __dut__._2509_/A __dut__._2863_/Q VGND VGND VPWR VPWR __dut__._1587_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2208_ __dut__._2208_/A1 __dut__._2208_/A2 __dut__._2207_/X VGND VGND VPWR
+ VPWR __dut__._2208_/X sky130_fd_sc_hd__a21o_4
XANTENNA__266__CLK _274_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2139_ __dut__._2141_/A __dut__._2139_/B VGND VGND VPWR VPWR __dut__._2139_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_146_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2992__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1971__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_168_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1960_ __dut__.__uuf__._1960_/A VGND VGND VPWR VPWR __dut__.__uuf__._1960_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1891_ __dut__.__uuf__._1923_/A __dut__.__uuf__._1891_/B __dut__.__uuf__._1891_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1892_/A sky130_fd_sc_hd__or3_4
XFILLER_149_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2307__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_11 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2032_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_136_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_22 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2010_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_117_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_33 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2138_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_55 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2318_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_44 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2224_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_155_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_77 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1398_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_88 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2264_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_99 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1606_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_66 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1554_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_105_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1325_ __dut__.__uuf__._1335_/A VGND VGND VPWR VPWR __dut__.__uuf__._1325_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_120_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2490_ __dut__._2502_/A1 __dut__._2490_/A2 __dut__._2489_/X VGND VGND VPWR
+ VPWR __dut__._2490_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1256_ __dut__._2369_/B __dut__.__uuf__._1025_/X __dut__.__uuf__._1219_/B
+ __dut__.__uuf__._1255_/X VGND VGND VPWR VPWR __dut__._2368_/A2 sky130_fd_sc_hd__o22a_4
X__dut__._1510_ __dut__._1510_/A1 __dut__._1508_/X __dut__._1509_/X VGND VGND VPWR
+ VPWR __dut__._2843_/D sky130_fd_sc_hd__a21o_4
XFILLER_74_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1441_ __dut__._1441_/A __dut__._2825_/Q VGND VGND VPWR VPWR __dut__._1441_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1187_ __dut__.__uuf__._1191_/A VGND VGND VPWR VPWR __dut__.__uuf__._1187_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1372_ rst VGND VGND VPWR VPWR __dut__._1372_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__289__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1018__A __dut__.__uuf__._1549_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1996__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._3042_ _271_/CLK __dut__._3042_/D __dut__._2576_/Y VGND VGND VPWR VPWR __dut__._3042_/Q
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._3023__D __dut__._3023_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2865__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_251_ _198_/X _251_/D VGND VGND VPWR VPWR _251_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_psn_inst_psn_buff_21_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_182_ _270_/Q _182_/B VGND VGND VPWR VPWR _269_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2217__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2826_ __dut__._2836_/CLK __dut__._2826_/D __dut__._2792_/Y VGND VGND VPWR
+ VPWR __dut__._2826_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2757_ rst VGND VGND VPWR VPWR __dut__._2757_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1708_ __dut__._1714_/A1 tie[6] __dut__._1707_/X VGND VGND VPWR VPWR __dut__._2911_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_2_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2688_ rst VGND VGND VPWR VPWR __dut__._2688_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1639_ __dut__._2457_/A __dut__._2876_/Q VGND VGND VPWR VPWR __dut__._1639_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3020__CLK clkbuf_opt_2_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_285_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2164__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1110_ __dut__.__uuf__._1117_/A VGND VGND VPWR VPWR __dut__.__uuf__._1110_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2090_ VGND VGND VPWR VPWR __dut__.__uuf__._2090_/HI tie[97] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2797__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1041_ __dut__.__uuf__._1019_/X __dut__.__uuf__._1040_/X prod[59]
+ prod[60] __dut__.__uuf__._1036_/X VGND VGND VPWR VPWR __dut__._2500_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._2888__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1978__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1943_ __dut__.__uuf__._1943_/A VGND VGND VPWR VPWR __dut__.__uuf__._1945_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1874_ __dut__._2195_/B __dut__._2201_/B VGND VGND VPWR VPWR __dut__.__uuf__._1875_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_149_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1990_ __dut__._1990_/A1 tie[147] __dut__._1989_/X VGND VGND VPWR VPWR __dut__._3052_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_137_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1902__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1565__A2 __dut__.__uuf__._1828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2611_ rst VGND VGND VPWR VPWR __dut__._2611_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2357_ __dut__.__uuf__._2358_/CLK __dut__._2494_/X __dut__.__uuf__._1048_/X
+ VGND VGND VPWR VPWR prod[56] sky130_fd_sc_hd__dfrtp_4
XFILLER_120_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2542_ rst VGND VGND VPWR VPWR __dut__._2542_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._1020__B __dut__._2109_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2288_ __dut__.__uuf__._2288_/CLK __dut__._2356_/X __dut__.__uuf__._1286_/X
+ VGND VGND VPWR VPWR __dut__._2357_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1308_ __dut__.__uuf__._1308_/A VGND VGND VPWR VPWR __dut__.__uuf__._1308_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1239_ __dut__.__uuf__._1254_/A VGND VGND VPWR VPWR __dut__.__uuf__._1239_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_115_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2473_ __dut__._2491_/A prod[45] VGND VGND VPWR VPWR __dut__._2473_/X sky130_fd_sc_hd__and2_4
XFILLER_74_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1424_ __dut__._1374_/Y mc[20] __dut__._1423_/X VGND VGND VPWR VPWR __dut__._1424_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_28_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_69_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_tck clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR clkbuf_3_3_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_131_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3025_ clkbuf_5_0_0_tck/X __dut__._3025_/D __dut__._2593_/Y VGND VGND VPWR
+ VPWR __dut__._3025_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._3043__CLK __dut__._3058_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_303_ _315_/CLK _303_/D trst VGND VGND VPWR VPWR _303_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_234_ _234_/A _234_/B VGND VGND VPWR VPWR _305_/D sky130_fd_sc_hd__and2_4
XFILLER_24_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2394__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_165_ _183_/A VGND VGND VPWR VPWR _173_/B sky130_fd_sc_hd__buf_2
XFILLER_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2809_ rst VGND VGND VPWR VPWR __dut__._2809_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1590_ __dut__.__uuf__._1590_/A VGND VGND VPWR VPWR __dut__.__uuf__._1590_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2211_ __dut__.__uuf__._2230_/CLK __dut__._2202_/X __dut__.__uuf__._1588_/X
+ VGND VGND VPWR VPWR __dut__._2203_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2142_ VGND VGND VPWR VPWR __dut__.__uuf__._2142_/HI tie[149] sky130_fd_sc_hd__conb_1
XFILLER_142_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2073_ VGND VGND VPWR VPWR __dut__.__uuf__._2073_/HI tie[80] sky130_fd_sc_hd__conb_1
XFILLER_29_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1024_ __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR __dut__.__uuf__._1229_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_96_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3066__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_209 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1963_/A sky130_fd_sc_hd__buf_2
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1926_ __dut__.__uuf__._1926_/A VGND VGND VPWR VPWR __dut__.__uuf__._1975_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_61_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1857_ __dut__.__uuf__._1813_/X __dut__.__uuf__._1855_/B __dut__.__uuf__._1855_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1858_/C sky130_fd_sc_hd__o21a_4
XANTENNA___dut__.__uuf__._2196__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1788_ __dut__.__uuf__._1788_/A VGND VGND VPWR VPWR __dut__.__uuf__._1788_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_137_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1973_ __dut__._2005_/A __dut__._3043_/Q VGND VGND VPWR VPWR __dut__._1973_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_3_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2525_ rst VGND VGND VPWR VPWR __dut__._2525_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2456_ __dut__._2502_/A1 __dut__._2456_/A2 __dut__._2455_/X VGND VGND VPWR
+ VPWR __dut__._2456_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1407_ __dut__._2509_/A __dut__._2818_/Q VGND VGND VPWR VPWR __dut__._1407_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2387_ __dut__._2389_/A prod[2] VGND VGND VPWR VPWR __dut__._2387_/X sky130_fd_sc_hd__and2_4
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3008_ _274_/CLK __dut__._3008_/D __dut__._2610_/Y VGND VGND VPWR VPWR __dut__._3008_/Q
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1206__A __dut__.__uuf__._1463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_217_ _293_/Q _232_/A VGND VGND VPWR VPWR _292_/D sky130_fd_sc_hd__and2_4
XFILLER_144_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_148_ _309_/Q _146_/Y _296_/Q _147_/X VGND VGND VPWR VPWR _309_/D sky130_fd_sc_hd__a211o_4
XANTENNA___dut__._2405__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_opt_2_tck_A clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3089__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_248_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_150_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1711_ __dut__._1596_/X VGND VGND VPWR VPWR __dut__.__uuf__._1715_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2926__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0___dut__.__uuf__.__clk_source__ clkbuf_2_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._2358__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1642_ __dut__.__uuf__._1645_/A VGND VGND VPWR VPWR __dut__.__uuf__._1642_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1573_ __dut__.__uuf__._1597_/A VGND VGND VPWR VPWR __dut__.__uuf__._1578_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2315__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2125_ VGND VGND VPWR VPWR __dut__.__uuf__._2125_/HI tie[132] sky130_fd_sc_hd__conb_1
XFILLER_102_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._2056_ VGND VGND VPWR VPWR __dut__.__uuf__._2056_/HI tie[63] sky130_fd_sc_hd__conb_1
X__dut__._2310_ __dut__._2310_/A1 __dut__._2310_/A2 __dut__._2309_/X VGND VGND VPWR
+ VPWR __dut__._2310_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2241_ __dut__._2245_/A __dut__._2241_/B VGND VGND VPWR VPWR __dut__._2241_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_112_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2172_ __dut__._2172_/A1 __dut__._2172_/A2 __dut__._2171_/X VGND VGND VPWR
+ VPWR __dut__._2172_/X sky130_fd_sc_hd__a21o_4
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1909_ __dut__.__uuf__._1952_/A __dut__.__uuf__._1909_/B __dut__.__uuf__._1909_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1910_/A sky130_fd_sc_hd__or3_4
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2225__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1956_ __dut__._1956_/A1 tie[130] __dut__._1955_/X VGND VGND VPWR VPWR __dut__._3035_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1572__A2 mp[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1887_ __dut__._2081_/A __dut__._3000_/Q VGND VGND VPWR VPWR __dut__._1887_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__.__uuf__._2211__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_121_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2508_ __dut__._2508_/A1 __dut__._2508_/A2 __dut__._2507_/X VGND VGND VPWR
+ VPWR __dut__._2508_/X sky130_fd_sc_hd__a21o_4
XFILLER_75_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2439_ __dut__._2507_/A prod[28] VGND VGND VPWR VPWR __dut__._2439_/X sky130_fd_sc_hd__and2_4
XFILLER_90_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3104__CLK __dut__._3106_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1625_ __dut__.__uuf__._1627_/A VGND VGND VPWR VPWR __dut__.__uuf__._1625_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2045__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1810_ __dut__._1816_/A1 tie[57] __dut__._1809_/X VGND VGND VPWR VPWR __dut__._2962_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1556_ __dut__.__uuf__._1562_/A VGND VGND VPWR VPWR __dut__.__uuf__._1556_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_123_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2234__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2790_ rst VGND VGND VPWR VPWR __dut__._2790_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1741_ __dut__._2189_/A __dut__._2927_/Q VGND VGND VPWR VPWR __dut__._1741_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1487_ __dut__.__uuf__._1550_/A VGND VGND VPWR VPWR __dut__.__uuf__._1487_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1672_ __dut__._2488_/A1 prod[53] __dut__._1671_/X VGND VGND VPWR VPWR __dut__._2893_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2108_ VGND VGND VPWR VPWR __dut__.__uuf__._2108_/HI tie[115] sky130_fd_sc_hd__conb_1
XFILLER_76_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2039_ VGND VGND VPWR VPWR __dut__.__uuf__._2039_/HI tie[46] sky130_fd_sc_hd__conb_1
XFILLER_123_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2224_ __dut__._2224_/A1 __dut__._2224_/A2 __dut__._2223_/X VGND VGND VPWR
+ VPWR __dut__._2224_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2155_ __dut__._2207_/A __dut__._2155_/B VGND VGND VPWR VPWR __dut__._2155_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_32_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2086_ __dut__._2488_/A1 prod[25] __dut__._2085_/X VGND VGND VPWR VPWR __dut__._3100_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2988_ __dut__._3096_/CLK __dut__._2988_/D __dut__._2630_/Y VGND VGND VPWR
+ VPWR __dut__._2988_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1939_ __dut__._2189_/A __dut__._3026_/Q VGND VGND VPWR VPWR __dut__._1939_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_113_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__292__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1536__A2 mp[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1410_ __dut__.__uuf__._1403_/X __dut__.__uuf__._1409_/X __dut__._2311_/B
+ __dut__.__uuf__._1403_/X VGND VGND VPWR VPWR __dut__._2310_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1341_ __dut__.__uuf__._1360_/A VGND VGND VPWR VPWR __dut__.__uuf__._1341_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_144_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1272_ __dut__.__uuf__._1292_/A VGND VGND VPWR VPWR __dut__.__uuf__._1492_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1472__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_5 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1924_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__309__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2911_ clkbuf_5_2_0_tck/X __dut__._2911_/D __dut__._2707_/Y VGND VGND VPWR
+ VPWR __dut__._2911_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1608_ __dut__.__uuf__._1609_/A VGND VGND VPWR VPWR __dut__.__uuf__._1608_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2842_ __dut__._2509_/B __dut__._2842_/D __dut__._2776_/Y VGND VGND VPWR
+ VPWR __dut__._2842_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1539_ __dut__.__uuf__._1528_/X __dut__.__uuf__._1523_/X __dut__._2253_/B
+ __dut__.__uuf__._1533_/X __dut__.__uuf__._1538_/X VGND VGND VPWR VPWR __dut__._2252_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._2773_ rst VGND VGND VPWR VPWR __dut__._2773_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1724_ __dut__._1726_/A1 tie[14] __dut__._1723_/X VGND VGND VPWR VPWR __dut__._2919_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_99_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1655_ __dut__._2491_/A __dut__._2884_/Q VGND VGND VPWR VPWR __dut__._1655_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1586_ __dut__._1780_/A1 __dut__._1584_/X __dut__._1585_/X VGND VGND VPWR
+ VPWR __dut__._2862_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_5_7_0_tck clkbuf_5_7_0_tck/A VGND VGND VPWR VPWR clkbuf_opt_2_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_94_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2207_ __dut__._2207_/A __dut__._2207_/B VGND VGND VPWR VPWR __dut__._2207_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2138_ __dut__._2138_/A1 __dut__._2138_/A2 __dut__._2137_/X VGND VGND VPWR
+ VPWR __dut__._2138_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2069_ __dut__._2069_/A __dut__._3091_/Q VGND VGND VPWR VPWR __dut__._2069_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1214__A __dut__.__uuf__._1214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_230_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1890_ __dut__.__uuf__._1867_/X __dut__.__uuf__._1888_/B __dut__.__uuf__._1888_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1891_/C sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._1699__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_12 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2030_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_136_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_23 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2008_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_34 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2140_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_56 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2368_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_45 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR psn_inst_psn_buff_57/A
+ sky130_fd_sc_hd__buf_2
XFILLER_145_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2323__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_78 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1714_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_89 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2266_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_67 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1598_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_132_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1324_ __dut__.__uuf__._1311_/X __dut__.__uuf__._1323_/X __dut__._2345_/B
+ __dut__.__uuf__._1311_/X VGND VGND VPWR VPWR __dut__._2344_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1255_ __dut__.__uuf__._1414_/A VGND VGND VPWR VPWR __dut__.__uuf__._1255_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1440_ __dut__._1374_/Y mc[24] __dut__._1439_/X VGND VGND VPWR VPWR __dut__._1440_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1186_ __dut__.__uuf__._1177_/X __dut__.__uuf__._1173_/X prod[10]
+ prod[11] __dut__.__uuf__._1185_/X VGND VGND VPWR VPWR __dut__._2402_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_104_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3041_ _315_/CLK __dut__._3041_/D __dut__._2577_/Y VGND VGND VPWR VPWR __dut__._3041_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_54_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_250_ _199_/X _314_/Q VGND VGND VPWR VPWR _250_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_181_ _271_/Q _182_/B VGND VGND VPWR VPWR _270_/D sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_14_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2825_ __dut__._2846_/CLK __dut__._2825_/D __dut__._2793_/Y VGND VGND VPWR
+ VPWR __dut__._2825_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2233__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2756_ rst VGND VGND VPWR VPWR __dut__._2756_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1707_ __dut__._2189_/A __dut__._2910_/Q VGND VGND VPWR VPWR __dut__._1707_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2687_ rst VGND VGND VPWR VPWR __dut__._2687_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1638_ __dut__._1638_/A1 prod[36] __dut__._1637_/X VGND VGND VPWR VPWR __dut__._2876_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1684__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1569_ __dut__._1569_/A __dut__._2857_/Q VGND VGND VPWR VPWR __dut__._1569_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_18_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1436__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0___dut__.__uuf__.__clk_source__ clkbuf_4_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2230_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2143__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_278_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1040_ __dut__.__uuf__._1099_/A VGND VGND VPWR VPWR __dut__.__uuf__._1040_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_83_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1942_ __dut__.__uuf__._1952_/A __dut__.__uuf__._1942_/B __dut__.__uuf__._1942_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1943_/A sky130_fd_sc_hd__or3_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1873_ __dut__._1424_/X VGND VGND VPWR VPWR __dut__.__uuf__._1877_/B
+ sky130_fd_sc_hd__inv_2
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._2053__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2610_ rst VGND VGND VPWR VPWR __dut__._2610_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1565__A3 __dut__._2239_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2356_ __dut__.__uuf__._2358_/CLK __dut__._2492_/X __dut__.__uuf__._1050_/X
+ VGND VGND VPWR VPWR prod[55] sky130_fd_sc_hd__dfrtp_4
XFILLER_105_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2541_ rst VGND VGND VPWR VPWR __dut__._2541_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2287_ __dut__.__uuf__._2307_/CLK __dut__._2354_/X __dut__.__uuf__._1290_/X
+ VGND VGND VPWR VPWR __dut__._2355_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1307_ __dut__.__uuf__._1300_/X __dut__.__uuf__._1306_/X __dut__._2351_/B
+ __dut__.__uuf__._1300_/X VGND VGND VPWR VPWR __dut__._2350_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1666__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2472_ __dut__._2488_/A1 __dut__._2472_/A2 __dut__._2471_/X VGND VGND VPWR
+ VPWR __dut__._2472_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1238_ __dut__.__uuf__._1340_/A VGND VGND VPWR VPWR __dut__.__uuf__._1254_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_101_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1423_ __dut__._2509_/A __dut__._2822_/Q VGND VGND VPWR VPWR __dut__._1423_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1169_ __dut__.__uuf__._1175_/A VGND VGND VPWR VPWR __dut__.__uuf__._1169_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2832__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1418__A1 __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3024_ clkbuf_5_1_0_tck/X __dut__._3024_/D __dut__._2594_/Y VGND VGND VPWR
+ VPWR __dut__._3024_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ _313_/CLK _302_/D trst VGND VGND VPWR VPWR _302_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_233_ _291_/Q _298_/Q _305_/Q _306_/Q VGND VGND VPWR VPWR _234_/B sky130_fd_sc_hd__or4_4
XFILLER_11_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_164_ _285_/Q _164_/B VGND VGND VPWR VPWR _284_/D sky130_fd_sc_hd__and2_4
XFILLER_136_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2808_ rst VGND VGND VPWR VPWR __dut__._2808_/Y sky130_fd_sc_hd__inv_2
X__dut__._2739_ rst VGND VGND VPWR VPWR __dut__._2739_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1977__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2210_ __dut__.__uuf__._2230_/CLK __dut__._2200_/X __dut__.__uuf__._1589_/X
+ VGND VGND VPWR VPWR __dut__._2201_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_154_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1896__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2601__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2141_ VGND VGND VPWR VPWR __dut__.__uuf__._2141_/HI tie[148] sky130_fd_sc_hd__conb_1
XFILLER_115_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._2855__CLK __dut__._2860_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2072_ VGND VGND VPWR VPWR __dut__.__uuf__._2072_/HI tie[79] sky130_fd_sc_hd__conb_1
XFILLER_68_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1648__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1023_ __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR __dut__.__uuf__._1023_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_45_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1925_ __dut__.__uuf__._1917_/A __dut__.__uuf__._1923_/B __dut__.__uuf__._1882_/X
+ VGND VGND VPWR VPWR __dut__._2210_/A2 sky130_fd_sc_hd__o21a_4
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1856_ __dut__.__uuf__._1856_/A VGND VGND VPWR VPWR __dut__.__uuf__._1858_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1787_ __dut__._2163_/B __dut__._2169_/B VGND VGND VPWR VPWR __dut__.__uuf__._1788_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_137_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1972_ __dut__._2004_/A1 tie[138] __dut__._1971_/X VGND VGND VPWR VPWR __dut__._3043_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_152_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2339_ __dut__.__uuf__._2358_/CLK __dut__._2458_/X __dut__.__uuf__._1101_/X
+ VGND VGND VPWR VPWR prod[38] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2511__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2524_ rst VGND VGND VPWR VPWR __dut__._2524_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_81_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2455_ __dut__._2457_/A prod[36] VGND VGND VPWR VPWR __dut__._2455_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1982__A __dut__.__uuf__._1982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3010__CLK _274_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1406_ __dut__._1418_/A1 __dut__._1404_/X __dut__._1405_/X VGND VGND VPWR
+ VPWR __dut__._2817_/D sky130_fd_sc_hd__a21o_4
X__dut__._2386_ __dut__._2412_/A1 __dut__._2386_/A2 __dut__._2385_/X VGND VGND VPWR
+ VPWR __dut__._2386_/X sky130_fd_sc_hd__a21o_4
XFILLER_74_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2064__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3007_ _274_/CLK __dut__._3007_/D __dut__._2611_/Y VGND VGND VPWR VPWR __dut__._3007_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_216_ _294_/Q _292_/Q _232_/A VGND VGND VPWR VPWR _291_/D sky130_fd_sc_hd__o21a_4
X_147_ _310_/Q _239_/A VGND VGND VPWR VPWR _147_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2405__B prod[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2290__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_144_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2878__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2421__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_143_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1710_ __dut__.__uuf__._1926_/A VGND VGND VPWR VPWR __dut__.__uuf__._1761_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1641_ __dut__.__uuf__._1645_/A VGND VGND VPWR VPWR __dut__.__uuf__._1641_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_119_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1572_ __dut__.__uuf__._1603_/A VGND VGND VPWR VPWR __dut__.__uuf__._1597_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_134_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_tck clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR clkbuf_3_1_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_143_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2124_ VGND VGND VPWR VPWR __dut__.__uuf__._2124_/HI tie[131] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._3033__CLK clkbuf_5_1_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2331__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2055_ VGND VGND VPWR VPWR __dut__.__uuf__._2055_/HI tie[62] sky130_fd_sc_hd__conb_1
XFILLER_110_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2240_ __dut__._2246_/A1 __dut__._2240_/A2 __dut__._2239_/X VGND VGND VPWR
+ VPWR __dut__._2240_/X sky130_fd_sc_hd__a21o_4
XFILLER_29_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2163__CLK __dut__.__uuf__._2303_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_112_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2046__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2171_ __dut__._2189_/A __dut__._2171_/B VGND VGND VPWR VPWR __dut__._2171_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1908_ __dut__._2207_/B __dut__._2213_/B __dut__.__uuf__._1907_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1909_/C sky130_fd_sc_hd__o21ai_4
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1839_ __dut__.__uuf__._1832_/A __dut__.__uuf__._1837_/B __dut__.__uuf__._1828_/X
+ VGND VGND VPWR VPWR __dut__._2178_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_40_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1955_ __dut__._2207_/A __dut__._3034_/Q VGND VGND VPWR VPWR __dut__._1955_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_137_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1886_ __dut__._1886_/A1 tie[95] __dut__._1885_/X VGND VGND VPWR VPWR __dut__._3000_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2507_ __dut__._2507_/A prod[62] VGND VGND VPWR VPWR __dut__._2507_/X sky130_fd_sc_hd__and2_4
X__dut__._2438_ __dut__._2438_/A1 __dut__._2438_/A2 __dut__._2437_/X VGND VGND VPWR
+ VPWR __dut__._2438_/X sky130_fd_sc_hd__a21o_4
XFILLER_75_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2369_ __dut__._2407_/A __dut__._2369_/B VGND VGND VPWR VPWR __dut__._2369_/X
+ sky130_fd_sc_hd__and2_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3056__CLK __dut__._3059_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2151__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_260_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__.__uuf__._2186__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_39_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1624_ __dut__.__uuf__._1627_/A VGND VGND VPWR VPWR __dut__.__uuf__._1624_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1555_ __dut__.__uuf__._1549_/X __dut__.__uuf__._1544_/X __dut__._2245_/B
+ __dut__.__uuf__._1447_/A __dut__.__uuf__._1554_/X VGND VGND VPWR VPWR __dut__._2244_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1740_ __dut__._1942_/A1 tie[22] __dut__._1739_/X VGND VGND VPWR VPWR __dut__._2927_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1486_ __dut__.__uuf__._1549_/A VGND VGND VPWR VPWR __dut__.__uuf__._1486_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1671_ __dut__._2491_/A __dut__._2892_/Q VGND VGND VPWR VPWR __dut__._1671_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2061__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2107_ VGND VGND VPWR VPWR __dut__.__uuf__._2107_/HI tie[114] sky130_fd_sc_hd__conb_1
XFILLER_130_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_opt_0_tck clkbuf_opt_2_tck/A VGND VGND VPWR VPWR clkbuf_opt_0_tck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2038_ VGND VGND VPWR VPWR __dut__.__uuf__._2038_/HI tie[45] sky130_fd_sc_hd__conb_1
XFILLER_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1405__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2223_ __dut__._2325_/A __dut__._2223_/B VGND VGND VPWR VPWR __dut__._2223_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2154_ __dut__._2172_/A1 __dut__._2154_/A2 __dut__._2153_/X VGND VGND VPWR
+ VPWR __dut__._2154_/X sky130_fd_sc_hd__a21o_4
XFILLER_53_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_44_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_opt_1_tck_A clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2085_ __dut__._2431_/A __dut__._3099_/Q VGND VGND VPWR VPWR __dut__._2085_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2987_ __dut__._3096_/CLK __dut__._2987_/D __dut__._2631_/Y VGND VGND VPWR
+ VPWR __dut__._2987_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1938_ __dut__._1942_/A1 tie[121] __dut__._1937_/X VGND VGND VPWR VPWR __dut__._3026_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1869_ __dut__._1881_/A __dut__._2991_/Q VGND VGND VPWR VPWR __dut__._1869_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2916__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_106_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1985__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1340_ __dut__.__uuf__._1340_/A VGND VGND VPWR VPWR __dut__.__uuf__._1360_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_113_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1271_ __dut__.__uuf__._1311_/A VGND VGND VPWR VPWR __dut__.__uuf__._1271_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_112_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1472__A2 mc[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2201__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_6 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1922_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2910_ clkbuf_5_2_0_tck/X __dut__._2910_/D __dut__._2708_/Y VGND VGND VPWR
+ VPWR __dut__._2910_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1895__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1044__B1 prod[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1607_ __dut__.__uuf__._1609_/A VGND VGND VPWR VPWR __dut__.__uuf__._1607_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_118_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2841_ __dut__._2509_/B __dut__._2841_/D __dut__._2777_/Y VGND VGND VPWR
+ VPWR __dut__._2841_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2772_ rst VGND VGND VPWR VPWR __dut__._2772_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1538_ __dut__._1504_/X __dut__.__uuf__._1529_/X __dut__._2255_/B
+ __dut__.__uuf__._1534_/X VGND VGND VPWR VPWR __dut__.__uuf__._1538_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__.__uuf__._1320__A __dut__.__uuf__._1709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2503__B prod[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1723_ __dut__._2189_/A __dut__._2918_/Q VGND VGND VPWR VPWR __dut__._1723_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2488__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1469_ __dut__.__uuf__._1533_/A VGND VGND VPWR VPWR __dut__.__uuf__._1469_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1654_ __dut__._2488_/A1 prod[44] __dut__._1653_/X VGND VGND VPWR VPWR __dut__._2884_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._3037__D __dut__._3037_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1585_ __dut__._1589_/A __dut__._2861_/Q VGND VGND VPWR VPWR __dut__._1585_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2206_ __dut__._2208_/A1 __dut__._2206_/A2 __dut__._2205_/X VGND VGND VPWR
+ VPWR __dut__._2206_/X sky130_fd_sc_hd__a21o_4
X__dut__._2137_ __dut__._2141_/A __dut__._2137_/B VGND VGND VPWR VPWR __dut__._2137_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2412__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2068_ __dut__._2422_/A1 prod[16] __dut__._2067_/X VGND VGND VPWR VPWR __dut__._3091_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_139_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_223_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2224__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_91_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_190 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._2192_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_13 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2028_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_118_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1026__B1 __dut__._2113_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2604__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_24 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2006_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_35 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2134_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_46 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2232_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_79 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1410_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_68 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1438_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1140__A __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1041__A3 prod[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_57 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2120_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1323_ __dut__.__uuf__._1319_/Y __dut__.__uuf__._1321_/X __dut__.__uuf__._1322_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1323_/X sky130_fd_sc_hd__o21a_4
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1254_ __dut__.__uuf__._1254_/A VGND VGND VPWR VPWR __dut__.__uuf__._1254_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1185_ __dut__.__uuf__._1200_/A VGND VGND VPWR VPWR __dut__.__uuf__._1185_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_74_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._3040_ _306_/CLK __dut__._3040_/D __dut__._2578_/Y VGND VGND VPWR VPWR __dut__._3040_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_120_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_180_ _272_/Q _187_/B VGND VGND VPWR VPWR _271_/D sky130_fd_sc_hd__or2_4
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2514__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2824_ __dut__._2846_/CLK __dut__._2824_/D __dut__._2794_/Y VGND VGND VPWR
+ VPWR __dut__._2824_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2755_ rst VGND VGND VPWR VPWR __dut__._2755_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1706_ __dut__._1714_/A1 tie[5] __dut__._1705_/X VGND VGND VPWR VPWR __dut__._2910_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2686_ rst VGND VGND VPWR VPWR __dut__._2686_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1637_ __dut__._2507_/A __dut__._2875_/Q VGND VGND VPWR VPWR __dut__._1637_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1684__A2 prod[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1568_ __dut__._1374_/Y mp[21] __dut__._1567_/X VGND VGND VPWR VPWR __dut__._1568_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_92_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1499_ __dut__._2509_/A __dut__._2841_/Q VGND VGND VPWR VPWR __dut__._1499_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1436__A2 mc[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_173_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1941_ __dut__._2219_/B __dut__._2225_/B __dut__.__uuf__._1940_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1942_/C sky130_fd_sc_hd__o21ai_4
XANTENNA___dut__._1503__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1872_ __dut__.__uuf__._1926_/A VGND VGND VPWR VPWR __dut__.__uuf__._1923_/A
+ sky130_fd_sc_hd__buf_2
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_6_0_tck clkbuf_5_7_0_tck/A VGND VGND VPWR VPWR clkbuf_5_6_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2355_ __dut__.__uuf__._2358_/CLK __dut__._2490_/X __dut__.__uuf__._1053_/X
+ VGND VGND VPWR VPWR prod[54] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_4_11_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2358_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1306_ __dut__.__uuf__._1305_/Y __dut__.__uuf__._1294_/X __dut__.__uuf__._1296_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1306_/X sky130_fd_sc_hd__o21a_4
XFILLER_132_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2540_ rst VGND VGND VPWR VPWR __dut__._2540_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2286_ __dut__.__uuf__._2307_/CLK __dut__._2352_/X __dut__.__uuf__._1299_/X
+ VGND VGND VPWR VPWR __dut__._2353_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2471_ __dut__._2491_/A prod[44] VGND VGND VPWR VPWR __dut__._2471_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1237_ __dut__.__uuf__._1640_/A VGND VGND VPWR VPWR __dut__.__uuf__._1340_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1168_ __dut__.__uuf__._1162_/X __dut__.__uuf__._1159_/X prod[16]
+ prod[17] __dut__.__uuf__._1156_/X VGND VGND VPWR VPWR __dut__._2414_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1422_ __dut__._2288_/A1 __dut__._1420_/X __dut__._1421_/X VGND VGND VPWR
+ VPWR __dut__._2821_/D sky130_fd_sc_hd__a21o_4
XFILLER_101_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1099_ __dut__.__uuf__._1099_/A VGND VGND VPWR VPWR __dut__.__uuf__._1099_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2509__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3023_ clkbuf_5_3_0_tck/X __dut__._3023_/D __dut__._2595_/Y VGND VGND VPWR
+ VPWR __dut__._3023_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1413__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_301_ _313_/CLK _301_/D trst VGND VGND VPWR VPWR _301_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1045__A __dut__.__uuf__._1992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_232_ _232_/A _232_/B VGND VGND VPWR VPWR _304_/D sky130_fd_sc_hd__and2_4
XFILLER_156_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_163_ _286_/Q _172_/B VGND VGND VPWR VPWR _285_/D sky130_fd_sc_hd__or2_4
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2807_ rst VGND VGND VPWR VPWR __dut__._2807_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2738_ rst VGND VGND VPWR VPWR __dut__._2738_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2669_ rst VGND VGND VPWR VPWR __dut__._2669_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_290_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1993__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2140_ VGND VGND VPWR VPWR __dut__.__uuf__._2140_/HI tie[147] sky130_fd_sc_hd__conb_1
XFILLER_114_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2071_ VGND VGND VPWR VPWR __dut__.__uuf__._2071_/HI tie[78] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1022_ __dut__.__uuf__._1464_/A VGND VGND VPWR VPWR __dut__.__uuf__._1936_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2329__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1924_ __dut__.__uuf__._1924_/A VGND VGND VPWR VPWR __dut__._2212_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1855_ __dut__.__uuf__._1898_/A __dut__.__uuf__._1855_/B __dut__.__uuf__._1855_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1856_/A sky130_fd_sc_hd__or3_4
XFILLER_138_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1786_ __dut__._1388_/X VGND VGND VPWR VPWR __dut__.__uuf__._1790_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1584__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1971_ __dut__._2005_/A __dut__._3042_/Q VGND VGND VPWR VPWR __dut__._1971_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._2338_ __dut__.__uuf__._2364_/CLK __dut__._2456_/X __dut__.__uuf__._1106_/X
+ VGND VGND VPWR VPWR prod[37] sky130_fd_sc_hd__dfrtp_4
XFILLER_121_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2269_ __dut__.__uuf__._2278_/CLK __dut__._2318_/X __dut__.__uuf__._1386_/X
+ VGND VGND VPWR VPWR __dut__._2319_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2523_ rst VGND VGND VPWR VPWR __dut__._2523_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2454_ __dut__._2454_/A1 __dut__._2454_/A2 __dut__._2453_/X VGND VGND VPWR
+ VPWR __dut__._2454_/X sky130_fd_sc_hd__a21o_4
XFILLER_75_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1405_ __dut__._2189_/A __dut__._2816_/Q VGND VGND VPWR VPWR __dut__._1405_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_74_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2385_ __dut__._2385_/A prod[1] VGND VGND VPWR VPWR __dut__._2385_/X sky130_fd_sc_hd__and2_4
XFILLER_28_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3006_ _194_/A __dut__._3006_/D __dut__._2612_/Y VGND VGND VPWR VPWR __dut__._3006_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_70_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_215_ _225_/B VGND VGND VPWR VPWR _232_/A sky130_fd_sc_hd__buf_2
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_146_ _239_/A VGND VGND VPWR VPWR _146_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2702__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_136_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2149__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1640_ __dut__.__uuf__._1640_/A VGND VGND VPWR VPWR __dut__.__uuf__._1645_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1571_ __dut__.__uuf__._1571_/A VGND VGND VPWR VPWR __dut__.__uuf__._1571_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_119_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2822__CLK __dut__._2846_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2612__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2123_ VGND VGND VPWR VPWR __dut__.__uuf__._2123_/HI tie[130] sky130_fd_sc_hd__conb_1
XFILLER_69_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2054_ VGND VGND VPWR VPWR __dut__.__uuf__._2054_/HI tie[61] sky130_fd_sc_hd__conb_1
XFILLER_84_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2170_ __dut__._2172_/A1 __dut__._2170_/A2 __dut__._2169_/X VGND VGND VPWR
+ VPWR __dut__._2170_/X sky130_fd_sc_hd__a21o_4
XFILLER_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2059__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1907_ __dut__.__uuf__._1907_/A VGND VGND VPWR VPWR __dut__.__uuf__._1907_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1838_ __dut__.__uuf__._1838_/A VGND VGND VPWR VPWR __dut__._2180_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_138_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1769_ __dut__.__uuf__._1790_/A __dut__.__uuf__._1769_/B __dut__.__uuf__._1769_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1770_/A sky130_fd_sc_hd__or3_4
XFILLER_119_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1954_ __dut__._1954_/A1 tie[129] __dut__._1953_/X VGND VGND VPWR VPWR __dut__._3034_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_153_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2522__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1885_ __dut__._2081_/A __dut__._2999_/Q VGND VGND VPWR VPWR __dut__._1885_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2506_ __dut__._2506_/A1 __dut__._2506_/A2 __dut__._2505_/X VGND VGND VPWR
+ VPWR __dut__._2506_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_8_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2437_ __dut__._2507_/A prod[27] VGND VGND VPWR VPWR __dut__._2437_/X sky130_fd_sc_hd__and2_4
XFILLER_75_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2368_ __dut__._2368_/A1 __dut__._2368_/A2 __dut__._2367_/X VGND VGND VPWR
+ VPWR __dut__._2368_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__269__CLK _274_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_4_0___dut__.__uuf__.__clk_source___A clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2299_ __dut__._2303_/A __dut__._2299_/B VGND VGND VPWR VPWR __dut__._2299_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_31_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2845__CLK __dut__._2846_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1548__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._2995__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_129_ _121_/Y _231_/A _125_/X _128_/X VGND VGND VPWR VPWR _130_/A sky130_fd_sc_hd__a211o_4
XFILLER_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_253_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2607__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1511__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1623_ __dut__.__uuf__._1627_/A VGND VGND VPWR VPWR __dut__.__uuf__._1623_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1554_ __dut__._1488_/X __dut__.__uuf__._1550_/X __dut__._2247_/B
+ __dut__.__uuf__._1294_/A VGND VGND VPWR VPWR __dut__.__uuf__._1554_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1485_ __dut__.__uuf__._1501_/A VGND VGND VPWR VPWR __dut__.__uuf__._1485_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1670_ __dut__._2488_/A1 prod[52] __dut__._1669_/X VGND VGND VPWR VPWR __dut__._2892_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2106_ VGND VGND VPWR VPWR __dut__.__uuf__._2106_/HI tie[113] sky130_fd_sc_hd__conb_1
XFILLER_103_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2037_ VGND VGND VPWR VPWR __dut__.__uuf__._2037_/HI tie[44] sky130_fd_sc_hd__conb_1
XFILLER_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2222_ __dut__._2222_/A1 __dut__._2222_/A2 __dut__._2221_/X VGND VGND VPWR
+ VPWR __dut__._2222_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2153_ __dut__._2207_/A __dut__._2153_/B VGND VGND VPWR VPWR __dut__._2153_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_25_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2084_ __dut__._2488_/A1 prod[24] __dut__._2083_/X VGND VGND VPWR VPWR __dut__._3099_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_37_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2517__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1421__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1950__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2986_ __dut__._3096_/CLK __dut__._2986_/D __dut__._2632_/Y VGND VGND VPWR
+ VPWR __dut__._2986_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1937_ __dut__._2189_/A __dut__._3025_/Q VGND VGND VPWR VPWR __dut__._1937_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1868_ __dut__._1868_/A1 tie[86] __dut__._1867_/X VGND VGND VPWR VPWR __dut__._2991_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1799_ __dut__._2507_/A __dut__._2956_/Q VGND VGND VPWR VPWR __dut__._1799_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3023__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1270_ __dut__.__uuf__._1280_/A VGND VGND VPWR VPWR __dut__.__uuf__._1270_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2337__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_7 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1920_/A1 sky130_fd_sc_hd__buf_2
XFILLER_10_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2840_ __dut__._2509_/B __dut__._2840_/D __dut__._2778_/Y VGND VGND VPWR
+ VPWR __dut__._2840_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1606_ __dut__.__uuf__._1609_/A VGND VGND VPWR VPWR __dut__.__uuf__._1606_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1537_ __dut__.__uuf__._1543_/A VGND VGND VPWR VPWR __dut__.__uuf__._1537_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2771_ rst VGND VGND VPWR VPWR __dut__._2771_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1722_ __dut__._1760_/A1 tie[13] __dut__._1721_/X VGND VGND VPWR VPWR __dut__._2918_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1468_ __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR __dut__.__uuf__._1468_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_103_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2800__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1653_ __dut__._2491_/A __dut__._2883_/Q VGND VGND VPWR VPWR __dut__._1653_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1399_ __dut__.__uuf__._1399_/A VGND VGND VPWR VPWR __dut__.__uuf__._1399_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_134_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1584_ __dut__._1374_/Y mp[25] __dut__._1583_/X VGND VGND VPWR VPWR __dut__._1584_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_45_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2205_ __dut__._2207_/A __dut__._2205_/B VGND VGND VPWR VPWR __dut__._2205_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._3046__CLK __dut__._3058_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2136_ __dut__._2136_/A1 __dut__._2136_/A2 __dut__._2135_/X VGND VGND VPWR
+ VPWR __dut__._2136_/X sky130_fd_sc_hd__a21o_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2067_ __dut__._2415_/A __dut__._3090_/Q VGND VGND VPWR VPWR __dut__._2067_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2969_ __dut__._2985_/CLK __dut__._2969_/D __dut__._2649_/Y VGND VGND VPWR
+ VPWR __dut__._2969_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2710__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_216_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2157__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_180 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._1626_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_191 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR psn_inst_psn_buff_201/A
+ sky130_fd_sc_hd__buf_2
XFILLER_31_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1026__B2 __dut__.__uuf__._1025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_14 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2026_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1914__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_25 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1960_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_36 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2136_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_47 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2234_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_69 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1434_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_58 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2230_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_132_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1322_ __dut__.__uuf__._1322_/A VGND VGND VPWR VPWR __dut__.__uuf__._1322_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1253_ __dut__.__uuf__._1248_/B __dut__.__uuf__._1251_/X __dut__.__uuf__._1214_/X
+ __dut__._2371_/B __dut__.__uuf__._1311_/A VGND VGND VPWR VPWR __dut__._2370_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_113_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2620__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_opt_0_tck_A clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1184_ __dut__.__uuf__._1191_/A VGND VGND VPWR VPWR __dut__.__uuf__._1184_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._3069__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__.__uuf__._2199__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2158__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2823_ __dut__._2846_/CLK __dut__._2823_/D __dut__._2795_/Y VGND VGND VPWR
+ VPWR __dut__._2823_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2754_ rst VGND VGND VPWR VPWR __dut__._2754_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1705_ __dut__._2189_/A __dut__._2909_/Q VGND VGND VPWR VPWR __dut__._1705_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_150_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2330__A1 __dut__._2332_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2685_ rst VGND VGND VPWR VPWR __dut__._2685_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2530__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1636_ __dut__._2104_/A1 prod[35] __dut__._1635_/X VGND VGND VPWR VPWR __dut__._2875_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1567_ __dut__._2509_/A __dut__._2858_/Q VGND VGND VPWR VPWR __dut__._1567_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1498_ __dut__._1498_/A1 __dut__._1496_/X __dut__._1497_/X VGND VGND VPWR
+ VPWR __dut__._2840_/D sky130_fd_sc_hd__a21o_4
XFILLER_73_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2119_ __dut__._2325_/A __dut__._2119_/B VGND VGND VPWR VPWR __dut__._2119_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._3099_ __dut__._3102_/CLK __dut__._3099_/D __dut__._2519_/Y VGND VGND VPWR
+ VPWR __dut__._3099_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2705__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_166_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1940_ __dut__.__uuf__._1940_/A VGND VGND VPWR VPWR __dut__.__uuf__._1940_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1871_ __dut__.__uuf__._1863_/A __dut__.__uuf__._1869_/B __dut__.__uuf__._1828_/X
+ VGND VGND VPWR VPWR __dut__._2190_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_51_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2388__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2615__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2354_ __dut__.__uuf__._2358_/CLK __dut__._2488_/X __dut__.__uuf__._1056_/X
+ VGND VGND VPWR VPWR prod[53] sky130_fd_sc_hd__dfrtp_4
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1305_ __dut__._2353_/B VGND VGND VPWR VPWR __dut__.__uuf__._1305_/Y
+ sky130_fd_sc_hd__inv_2
Xclkbuf_3_3_0___dut__.__uuf__.__clk_source__ clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_7_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_132_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2285_ __dut__.__uuf__._2307_/CLK __dut__._2350_/X __dut__.__uuf__._1304_/X
+ VGND VGND VPWR VPWR __dut__._2351_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_87_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2470_ __dut__._2488_/A1 __dut__._2470_/A2 __dut__._2469_/X VGND VGND VPWR
+ VPWR __dut__._2470_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1236_ __dut__.__uuf__._1214_/A __dut__.__uuf__._1235_/X __dut__.__uuf__._1226_/B
+ __dut__._2379_/B __dut__.__uuf__._1232_/X VGND VGND VPWR VPWR __dut__._2378_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__.__uuf__._1183__B1 prod[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1167_ __dut__.__uuf__._1175_/A VGND VGND VPWR VPWR __dut__.__uuf__._1167_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1421_ __dut__._2325_/A __dut__._2810_/Q VGND VGND VPWR VPWR __dut__._1421_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_101_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1098_ __dut__.__uuf__._1101_/A VGND VGND VPWR VPWR __dut__.__uuf__._1098_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3022_ clkbuf_opt_0_tck/X __dut__._3022_/D __dut__._2596_/Y VGND VGND VPWR
+ VPWR __dut__._3022_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_300_ _313_/CLK _300_/D trst VGND VGND VPWR VPWR _300_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_231_ _231_/A _298_/Q _305_/Q VGND VGND VPWR VPWR _232_/B sky130_fd_sc_hd__or3_4
XFILLER_11_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_162_ _287_/Q _164_/B VGND VGND VPWR VPWR _286_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2525__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2806_ rst VGND VGND VPWR VPWR __dut__._2806_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2214__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_151_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2737_ rst VGND VGND VPWR VPWR __dut__._2737_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2668_ rst VGND VGND VPWR VPWR __dut__._2668_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1619_ __dut__._2509_/A __dut__._2871_/Q VGND VGND VPWR VPWR __dut__._1619_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2599_ rst VGND VGND VPWR VPWR __dut__._2599_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_283_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2070_ VGND VGND VPWR VPWR __dut__.__uuf__._2070_/HI tie[77] sky130_fd_sc_hd__conb_1
XFILLER_84_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1021_ __dut__.__uuf__._1441_/A VGND VGND VPWR VPWR __dut__.__uuf__._1464_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_110_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1923_ __dut__.__uuf__._1923_/A __dut__.__uuf__._1923_/B __dut__.__uuf__._1923_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1924_/A sky130_fd_sc_hd__or3_4
XFILLER_37_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._3107__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1854_ __dut__._2187_/B __dut__._2193_/B __dut__.__uuf__._1853_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1855_/C sky130_fd_sc_hd__o21ai_4
XFILLER_138_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1785_ __dut__.__uuf__._1778_/A __dut__.__uuf__._1783_/B __dut__.__uuf__._1774_/X
+ VGND VGND VPWR VPWR __dut__._2158_/A2 sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._2345__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1970_ __dut__._2004_/A1 tie[137] __dut__._1969_/X VGND VGND VPWR VPWR __dut__._3042_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1584__A2 mp[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2237__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2337_ __dut__.__uuf__._2364_/CLK __dut__._2454_/X __dut__.__uuf__._1108_/X
+ VGND VGND VPWR VPWR prod[36] sky130_fd_sc_hd__dfrtp_4
XFILLER_114_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2522_ rst VGND VGND VPWR VPWR __dut__._2522_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2268_ __dut__.__uuf__._2278_/CLK __dut__._2316_/X __dut__.__uuf__._1392_/X
+ VGND VGND VPWR VPWR __dut__._2317_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_59_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1219_ __dut__.__uuf__._1219_/A __dut__.__uuf__._1219_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1248_/B sky130_fd_sc_hd__or2_4
XFILLER_142_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2199_ __dut__.__uuf__._2230_/CLK __dut__._2178_/X __dut__.__uuf__._1602_/X
+ VGND VGND VPWR VPWR __dut__._2179_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2453_ __dut__._2507_/A prod[35] VGND VGND VPWR VPWR __dut__._2453_/X sky130_fd_sc_hd__and2_4
XFILLER_75_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1404_ __dut__._1374_/Y mc[16] __dut__._1403_/X VGND VGND VPWR VPWR __dut__._1404_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._2384_ __dut__._2412_/A1 __dut__._2384_/A2 __dut__._2383_/X VGND VGND VPWR
+ VPWR __dut__._2384_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_67_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2239__B __dut__._2239_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3005_ _194_/A __dut__._3005_/D __dut__._2613_/Y VGND VGND VPWR VPWR __dut__._3005_/Q
+ sky130_fd_sc_hd__dfrtp_4
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ _234_/A _214_/B VGND VGND VPWR VPWR _225_/B sky130_fd_sc_hd__nor2_4
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_145_ _239_/A _142_/Y tdi _310_/Q _144_/Y VGND VGND VPWR VPWR _310_/D sky130_fd_sc_hd__a32o_4
XFILLER_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_5_0_tck clkbuf_5_5_0_tck/A VGND VGND VPWR VPWR clkbuf_5_5_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_129_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2165__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1570_ __dut__.__uuf__._1571_/A VGND VGND VPWR VPWR __dut__.__uuf__._1570_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2122_ VGND VGND VPWR VPWR __dut__.__uuf__._2122_/HI tie[129] sky130_fd_sc_hd__conb_1
XFILLER_130_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2053_ VGND VGND VPWR VPWR __dut__.__uuf__._2053_/HI tie[60] sky130_fd_sc_hd__conb_1
XFILLER_69_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1906_ __dut__._2207_/B __dut__._2213_/B VGND VGND VPWR VPWR __dut__.__uuf__._1907_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2075__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1837_ __dut__.__uuf__._1869_/A __dut__.__uuf__._1837_/B __dut__.__uuf__._1837_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1838_/A sky130_fd_sc_hd__or3_4
XANTENNA___dut__.__uuf__._1604__A __dut__.__uuf__._1628_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1768_ __dut__._2155_/B __dut__._2161_/B __dut__.__uuf__._1767_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1769_/C sky130_fd_sc_hd__o21ai_4
X__dut__._1953_ __dut__._2207_/A __dut__._3033_/Q VGND VGND VPWR VPWR __dut__._1953_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1699_ __dut__.__uuf__._1699_/A VGND VGND VPWR VPWR __dut__.__uuf__._1699_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2803__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1884_ __dut__._1884_/A1 tie[94] __dut__._1883_/X VGND VGND VPWR VPWR __dut__._2999_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_137_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1419__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2505_ __dut__._2505_/A prod[61] VGND VGND VPWR VPWR __dut__._2505_/X sky130_fd_sc_hd__and2_4
X__dut__._2436_ __dut__._2436_/A1 __dut__._2436_/A2 __dut__._2435_/X VGND VGND VPWR
+ VPWR __dut__._2436_/X sky130_fd_sc_hd__a21o_4
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2367_ __dut__._2407_/A __dut__._2367_/B VGND VGND VPWR VPWR __dut__._2367_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2298_ __dut__._2300_/A1 __dut__._2298_/A2 __dut__._2297_/X VGND VGND VPWR
+ VPWR __dut__._2298_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1548__A2 mp[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2713__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_128_ _214_/B VGND VGND VPWR VPWR _128_/X sky130_fd_sc_hd__buf_2
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_246_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1484__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1999__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1622_ __dut__.__uuf__._1628_/A VGND VGND VPWR VPWR __dut__.__uuf__._1627_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_147_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2623__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1553_ __dut__.__uuf__._1562_/A VGND VGND VPWR VPWR __dut__.__uuf__._1553_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1484_ __dut__.__uuf__._1566_/A VGND VGND VPWR VPWR __dut__.__uuf__._1501_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_131_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2105_ VGND VGND VPWR VPWR __dut__.__uuf__._2105_/HI tie[112] sky130_fd_sc_hd__conb_1
XFILLER_130_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2036_ VGND VGND VPWR VPWR __dut__.__uuf__._2036_/HI tie[43] sky130_fd_sc_hd__conb_1
X__dut__._2221_ __dut__._2325_/A __dut__._2221_/B VGND VGND VPWR VPWR __dut__._2221_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2152_ __dut__._2208_/A1 __dut__._2152_/A2 __dut__._2151_/X VGND VGND VPWR
+ VPWR __dut__._2152_/X sky130_fd_sc_hd__a21o_4
X__dut__._2083_ __dut__._2431_/A __dut__._3098_/Q VGND VGND VPWR VPWR __dut__._2083_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2985_ __dut__._2985_/CLK __dut__._2985_/D __dut__._2633_/Y VGND VGND VPWR
+ VPWR __dut__._2985_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2533__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1936_ __dut__._1942_/A1 tie[120] __dut__._1935_/X VGND VGND VPWR VPWR __dut__._3025_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_153_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1867_ __dut__._1881_/A __dut__._2990_/Q VGND VGND VPWR VPWR __dut__._1867_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1798_ __dut__._1830_/A1 tie[51] __dut__._1797_/X VGND VGND VPWR VPWR __dut__._2956_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2419_ __dut__._2419_/A prod[18] VGND VGND VPWR VPWR __dut__._2419_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2708__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2443__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2618__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_8 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1918_/A1 sky130_fd_sc_hd__buf_2
XFILLER_50_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1605_ __dut__.__uuf__._1609_/A VGND VGND VPWR VPWR __dut__.__uuf__._1605_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2353__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1536_ __dut__.__uuf__._1528_/X __dut__.__uuf__._1523_/X __dut__._2255_/B
+ __dut__.__uuf__._1533_/X __dut__.__uuf__._1535_/X VGND VGND VPWR VPWR __dut__._2254_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_151_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2770_ rst VGND VGND VPWR VPWR __dut__._2770_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1721_ __dut__._2189_/A __dut__._2917_/Q VGND VGND VPWR VPWR __dut__._1721_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1467_ __dut__.__uuf__._1463_/X __dut__.__uuf__._1458_/X __dut__._2287_/B
+ __dut__.__uuf__._1447_/X __dut__.__uuf__._1466_/X VGND VGND VPWR VPWR __dut__._2286_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_150_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1652_ __dut__._2488_/A1 prod[43] __dut__._1651_/X VGND VGND VPWR VPWR __dut__._2883_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1398_ __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR __dut__.__uuf__._1398_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_134_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1583_ __dut__._2509_/A __dut__._2862_/Q VGND VGND VPWR VPWR __dut__._1583_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_85_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1448__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2019_ VGND VGND VPWR VPWR __dut__.__uuf__._2019_/HI tie[26] sky130_fd_sc_hd__conb_1
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2204_ __dut__._2204_/A1 __dut__._2204_/A2 __dut__._2203_/X VGND VGND VPWR
+ VPWR __dut__._2204_/X sky130_fd_sc_hd__a21o_4
X__dut__._2135_ __dut__._2141_/A __dut__._2135_/B VGND VGND VPWR VPWR __dut__._2135_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2528__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2066_ __dut__._2412_/A1 prod[15] __dut__._2065_/X VGND VGND VPWR VPWR __dut__._3090_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1620__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2968_ __dut__._2985_/CLK __dut__._2968_/D __dut__._2650_/Y VGND VGND VPWR
+ VPWR __dut__._2968_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1919_ __dut__._2207_/A __dut__._3016_/Q VGND VGND VPWR VPWR __dut__._1919_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_5_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2899_ _306_/CLK __dut__._2899_/D __dut__._2719_/Y VGND VGND VPWR VPWR __dut__._2899_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_110_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1607__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2100__A2 prod[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_111_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_209_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_181 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._1630_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_170 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2412_/A1 sky130_fd_sc_hd__buf_8
XFILLER_145_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_192 psn_inst_psn_buff_201/A VGND VGND VPWR VPWR __dut__._1510_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1026__A2 __dut__.__uuf__._1023_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_15 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2024_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_129_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_26 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1958_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_37 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2130_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2173__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2270__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_59 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1458_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_48 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2236_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_117_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1321_ __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR __dut__.__uuf__._1321_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1252_ __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR __dut__.__uuf__._1311_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_113_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1678__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1183_ __dut__.__uuf__._1177_/X __dut__.__uuf__._1173_/X prod[11]
+ prod[12] __dut__.__uuf__._1170_/X VGND VGND VPWR VPWR __dut__._2404_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__.__uuf__._1149__A __dut__.__uuf__._1640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2822_ __dut__._2846_/CLK __dut__._2822_/D __dut__._2796_/Y VGND VGND VPWR
+ VPWR __dut__._2822_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_145_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1519_ __dut__.__uuf__._1522_/A VGND VGND VPWR VPWR __dut__.__uuf__._1519_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2753_ rst VGND VGND VPWR VPWR __dut__._2753_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1704_ __dut__._1714_/A1 tie[4] __dut__._1703_/X VGND VGND VPWR VPWR __dut__._2909_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_77_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2684_ rst VGND VGND VPWR VPWR __dut__._2684_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1427__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_97_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1059__A __dut__.__uuf__._1992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1635_ __dut__._2103_/A __dut__._3109_/Q VGND VGND VPWR VPWR __dut__._1635_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._3013__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1566_ __dut__._1566_/A1 __dut__._1564_/X __dut__._1565_/X VGND VGND VPWR
+ VPWR __dut__._2857_/D sky130_fd_sc_hd__a21o_4
XFILLER_57_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1497_ __dut__._2189_/A __dut__._2839_/Q VGND VGND VPWR VPWR __dut__._1497_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3098_ __dut__._3102_/CLK __dut__._3098_/D __dut__._2520_/Y VGND VGND VPWR
+ VPWR __dut__._3098_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1256__A2 __dut__.__uuf__._1025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2118_ __dut__._2120_/A1 __dut__._2118_/A2 __dut__._2117_/X VGND VGND VPWR
+ VPWR __dut__._2118_/X sky130_fd_sc_hd__a21o_4
XFILLER_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2049_ __dut__._2407_/A __dut__._3081_/Q VGND VGND VPWR VPWR __dut__._2049_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_127_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2721__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_159_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1870_ __dut__.__uuf__._1870_/A VGND VGND VPWR VPWR __dut__._2192_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_149_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2631__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2353_ __dut__.__uuf__._2353_/CLK __dut__._2486_/X __dut__.__uuf__._1060_/X
+ VGND VGND VPWR VPWR prod[52] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3036__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1304_ __dut__.__uuf__._1308_/A VGND VGND VPWR VPWR __dut__.__uuf__._1304_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2284_ __dut__.__uuf__._2288_/CLK __dut__._2348_/X __dut__.__uuf__._1308_/X
+ VGND VGND VPWR VPWR __dut__._2349_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_115_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1235_ __dut__._2379_/B __dut__.__uuf__._1240_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1235_/X sky130_fd_sc_hd__or2_4
XFILLER_140_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1166_ __dut__.__uuf__._1162_/X __dut__.__uuf__._1159_/X prod[17]
+ prod[18] __dut__.__uuf__._1156_/X VGND VGND VPWR VPWR __dut__._2416_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1420_ __dut__._1374_/Y mc[1] __dut__._1419_/X VGND VGND VPWR VPWR __dut__._1420_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2166__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1097_ __dut__.__uuf__._1088_/X __dut__.__uuf__._1085_/X prod[40]
+ prod[41] __dut__.__uuf__._1096_/X VGND VGND VPWR VPWR __dut__._2462_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3021_ clkbuf_opt_1_tck/X __dut__._3021_/D __dut__._2597_/Y VGND VGND VPWR
+ VPWR __dut__._3021_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_230_ _234_/A _304_/Q VGND VGND VPWR VPWR _303_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2806__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1999_ VGND VGND VPWR VPWR __dut__.__uuf__._1999_/HI tie[6] sky130_fd_sc_hd__conb_1
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_161_ _288_/Q _172_/B VGND VGND VPWR VPWR _287_/D sky130_fd_sc_hd__or2_4
XFILLER_155_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_12_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2000__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3059__D __dut__._3059_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2805_ rst VGND VGND VPWR VPWR __dut__._2805_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2541__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2736_ rst VGND VGND VPWR VPWR __dut__._2736_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2667_ rst VGND VGND VPWR VPWR __dut__._2667_/Y sky130_fd_sc_hd__inv_2
XANTENNA__302__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1618_ __dut__._2376_/A1 __dut__._1616_/X __dut__._1617_/X VGND VGND VPWR
+ VPWR __dut__._2870_/D sky130_fd_sc_hd__a21o_4
X__dut__._2598_ rst VGND VGND VPWR VPWR __dut__._2598_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1549_ __dut__._1557_/A __dut__._2852_/Q VGND VGND VPWR VPWR __dut__._1549_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_61_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2716__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3059__CLK __dut__._3059_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_276_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2189__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_122_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1020_ __dut__._2107_/B __dut__._2109_/B VGND VGND VPWR VPWR __dut__.__uuf__._1441_/A
+ sky130_fd_sc_hd__or2_4
XFILLER_110_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2058__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1922_ __dut__.__uuf__._1921_/X __dut__.__uuf__._1919_/B __dut__.__uuf__._1919_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1923_/C sky130_fd_sc_hd__o21a_4
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1853_ __dut__.__uuf__._1853_/A VGND VGND VPWR VPWR __dut__.__uuf__._1853_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2626__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1784_ __dut__.__uuf__._1784_/A VGND VGND VPWR VPWR __dut__._2160_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_138_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2361__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2336_ __dut__.__uuf__._2364_/CLK __dut__._2452_/X __dut__.__uuf__._1110_/X
+ VGND VGND VPWR VPWR prod[35] sky130_fd_sc_hd__dfrtp_4
XFILLER_126_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2521_ rst VGND VGND VPWR VPWR __dut__._2521_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2267_ __dut__.__uuf__._2278_/CLK __dut__._2314_/X __dut__.__uuf__._1396_/X
+ VGND VGND VPWR VPWR __dut__._2315_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2452_ __dut__._2452_/A1 __dut__._2452_/A2 __dut__._2451_/X VGND VGND VPWR
+ VPWR __dut__._2452_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1218_ __dut__._2369_/B VGND VGND VPWR VPWR __dut__.__uuf__._1219_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_87_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1705__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1403_ __dut__._2509_/A __dut__._2817_/Q VGND VGND VPWR VPWR __dut__._1403_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2198_ __dut__.__uuf__._2230_/CLK __dut__._2176_/X __dut__.__uuf__._1605_/X
+ VGND VGND VPWR VPWR __dut__._2177_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_142_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2383_ __dut__._2385_/A prod[0] VGND VGND VPWR VPWR __dut__._2383_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1149_ __dut__.__uuf__._1640_/A VGND VGND VPWR VPWR __dut__.__uuf__._1208_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_83_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3004_ _194_/A __dut__._3004_/D __dut__._2614_/Y VGND VGND VPWR VPWR __dut__._3004_/Q
+ sky130_fd_sc_hd__dfrtp_4
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2536__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ tms VGND VGND VPWR VPWR _234_/A sky130_fd_sc_hd__inv_2
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_144_ _220_/A VGND VGND VPWR VPWR _144_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2719_ rst VGND VGND VPWR VPWR __dut__._2719_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1615__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._2460__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__295__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2181__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2121_ VGND VGND VPWR VPWR __dut__.__uuf__._2121_/HI tie[128] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2052_ VGND VGND VPWR VPWR __dut__.__uuf__._2052_/HI tie[59] sky130_fd_sc_hd__conb_1
XFILLER_111_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1905_ __dut__._1436_/X VGND VGND VPWR VPWR __dut__.__uuf__._1909_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2204__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1836_ __dut__.__uuf__._1813_/X __dut__.__uuf__._1834_/B __dut__.__uuf__._1834_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1837_/C sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1767_ __dut__.__uuf__._1767_/A VGND VGND VPWR VPWR __dut__.__uuf__._1767_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_125_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1698_ __dut__._2131_/B __dut__._2137_/B VGND VGND VPWR VPWR __dut__.__uuf__._1699_/A
+ sky130_fd_sc_hd__and2_4
X__dut__._1952_ __dut__._1952_/A1 tie[128] __dut__._1951_/X VGND VGND VPWR VPWR __dut__._3033_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_119_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1883_ __dut__._2081_/A __dut__._2998_/Q VGND VGND VPWR VPWR __dut__._1883_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2319_ __dut__.__uuf__._2328_/CLK __dut__._2418_/X __dut__.__uuf__._1161_/X
+ VGND VGND VPWR VPWR prod[18] sky130_fd_sc_hd__dfrtp_4
XFILLER_88_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2504_ __dut__._2504_/A1 __dut__._2504_/A2 __dut__._2503_/X VGND VGND VPWR
+ VPWR __dut__._2504_/X sky130_fd_sc_hd__a21o_4
XFILLER_101_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2435_ __dut__._2435_/A prod[26] VGND VGND VPWR VPWR __dut__._2435_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1435__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2366_ __dut__._2368_/A1 __dut__._2366_/A2 __dut__._2365_/X VGND VGND VPWR
+ VPWR __dut__._2366_/X sky130_fd_sc_hd__a21o_4
XFILLER_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2297_ __dut__._2297_/A __dut__._2297_/B VGND VGND VPWR VPWR __dut__._2297_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_102_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_127_ tms _257_/D _258_/Q _127_/D VGND VGND VPWR VPWR _214_/B sky130_fd_sc_hd__and4_4
XFILLER_125_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2891__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_141_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1484__A2 mp[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2227__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_81_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_239_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1621_ __dut__.__uuf__._1621_/A VGND VGND VPWR VPWR __dut__.__uuf__._1621_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_107_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1552_ __dut__.__uuf__._1549_/X __dut__.__uuf__._1544_/X __dut__._2247_/B
+ __dut__.__uuf__._1533_/X __dut__.__uuf__._1551_/X VGND VGND VPWR VPWR __dut__._2246_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__.__uuf__._1440__A __dut__.__uuf__._1463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1483_ __dut__.__uuf__._1603_/A VGND VGND VPWR VPWR __dut__.__uuf__._1566_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_143_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2104_ VGND VGND VPWR VPWR __dut__.__uuf__._2104_/HI tie[111] sky130_fd_sc_hd__conb_1
XFILLER_131_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2035_ VGND VGND VPWR VPWR __dut__.__uuf__._2035_/HI tie[42] sky130_fd_sc_hd__conb_1
X__dut__._2220_ __dut__._2220_/A1 __dut__._2220_/A2 __dut__._2219_/X VGND VGND VPWR
+ VPWR __dut__._2220_/X sky130_fd_sc_hd__a21o_4
XFILLER_25_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2151_ __dut__._2207_/A __dut__._2151_/B VGND VGND VPWR VPWR __dut__._2151_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2082_ __dut__._2428_/A1 prod[23] __dut__._2081_/X VGND VGND VPWR VPWR __dut__._3098_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_16_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1047__B1 prod[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._1819_ __dut__._1400_/X VGND VGND VPWR VPWR __dut__.__uuf__._1823_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2984_ __dut__._2985_/CLK __dut__._2984_/D __dut__._2634_/Y VGND VGND VPWR
+ VPWR __dut__._2984_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1935_ __dut__._2189_/A __dut__._3024_/Q VGND VGND VPWR VPWR __dut__._1935_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_153_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_4_0_tck clkbuf_5_5_0_tck/A VGND VGND VPWR VPWR clkbuf_5_4_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1866_ __dut__._1866_/A1 tie[85] __dut__._1865_/X VGND VGND VPWR VPWR __dut__._2990_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_79_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1797_ __dut__._1797_/A __dut__._2955_/Q VGND VGND VPWR VPWR __dut__._1797_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2418_ __dut__._2422_/A1 __dut__._2418_/A2 __dut__._2417_/X VGND VGND VPWR
+ VPWR __dut__._2418_/X sky130_fd_sc_hd__a21o_4
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2349_ __dut__._2407_/A __dut__._2349_/B VGND VGND VPWR VPWR __dut__._2349_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2724__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2406__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1_0_tck_A clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1435__A __dut__.__uuf__._1480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_9 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1916_/A1 sky130_fd_sc_hd__buf_2
XFILLER_148_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2634__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1044__A3 prod[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1604_ __dut__.__uuf__._1628_/A VGND VGND VPWR VPWR __dut__.__uuf__._1609_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_147_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1535_ __dut__._1512_/X __dut__.__uuf__._1529_/X __dut__._2257_/B
+ __dut__.__uuf__._1534_/X VGND VGND VPWR VPWR __dut__.__uuf__._1535_/X sky130_fd_sc_hd__o22a_4
XFILLER_151_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1720_ __dut__._1760_/A1 tie[12] __dut__._1719_/X VGND VGND VPWR VPWR __dut__._2917_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._1201__B1 prod[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1466_ __dut__._1580_/X __dut__.__uuf__._1465_/X __dut__._2289_/B
+ __dut__.__uuf__._1448_/X VGND VGND VPWR VPWR __dut__.__uuf__._1466_/X sky130_fd_sc_hd__o22a_4
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1651_ __dut__._2491_/A __dut__._2882_/Q VGND VGND VPWR VPWR __dut__._1651_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1397_ __dut__._2317_/B VGND VGND VPWR VPWR __dut__.__uuf__._1397_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_89_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1582_ __dut__._1780_/A1 __dut__._1580_/X __dut__._1581_/X VGND VGND VPWR
+ VPWR __dut__._2861_/D sky130_fd_sc_hd__a21o_4
XFILLER_134_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2018_ VGND VGND VPWR VPWR __dut__.__uuf__._2018_/HI tie[25] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._1448__A2 mc[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2809__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1713__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2203_ __dut__._2507_/A __dut__._2203_/B VGND VGND VPWR VPWR __dut__._2203_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_60_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2134_ __dut__._2134_/A1 __dut__._2134_/A2 __dut__._2133_/X VGND VGND VPWR
+ VPWR __dut__._2134_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_42_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1620__A2 mc[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2065_ __dut__._2415_/A __dut__._3089_/Q VGND VGND VPWR VPWR __dut__._2065_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2544__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1384__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2967_ __dut__._2985_/CLK __dut__._2967_/D __dut__._2651_/Y VGND VGND VPWR
+ VPWR __dut__._2967_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1991__A1 done VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1918_ __dut__._1918_/A1 tie[111] __dut__._1917_/X VGND VGND VPWR VPWR __dut__._3016_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_141_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3092__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2898_ _306_/CLK __dut__._2898_/D __dut__._2720_/Y VGND VGND VPWR VPWR __dut__._2898_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_122_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1849_ __dut__._1881_/A __dut__._2981_/Q VGND VGND VPWR VPWR __dut__._1849_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_110_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2719__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1623__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpsn_inst_psn_buff_171 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2422_/A1 sky130_fd_sc_hd__buf_2
XANTENNA_psn_inst_psn_buff_104_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_182 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._1634_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_160 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2454_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_193 psn_inst_psn_buff_201/A VGND VGND VPWR VPWR __dut__._1450_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1026__A3 prod[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_16 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2022_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_27 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1956_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_38 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2132_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_133_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1320_ __dut__.__uuf__._1709_/A VGND VGND VPWR VPWR __dut__.__uuf__._1649_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_49 psn_inst_psn_buff_57/A VGND VGND VPWR VPWR __dut__._2110_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_144_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1251_ __dut__._2371_/B __dut__._2369_/B VGND VGND VPWR VPWR __dut__.__uuf__._1251_/X
+ sky130_fd_sc_hd__or2_4
XFILLER_140_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1678__A2 prod[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1182_ __dut__.__uuf__._1191_/A VGND VGND VPWR VPWR __dut__.__uuf__._1182_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_113_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2629__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2821_ __dut__._2860_/CLK __dut__._2821_/D __dut__._2797_/Y VGND VGND VPWR
+ VPWR __dut__._2821_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1518_ __dut__.__uuf__._1507_/X __dut__.__uuf__._1502_/X __dut__._2263_/B
+ __dut__.__uuf__._1512_/X __dut__.__uuf__._1517_/X VGND VGND VPWR VPWR __dut__._2262_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._2752_ rst VGND VGND VPWR VPWR __dut__._2752_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1703_ __dut__._2189_/A __dut__._2908_/Q VGND VGND VPWR VPWR __dut__._1703_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1449_ __dut__._1600_/X __dut__.__uuf__._1442_/X __dut__._2297_/B
+ __dut__.__uuf__._1448_/X VGND VGND VPWR VPWR __dut__.__uuf__._1449_/X sky130_fd_sc_hd__o22a_4
X__dut__._2683_ rst VGND VGND VPWR VPWR __dut__._2683_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1634_ __dut__._1634_/A1 __dut__._1632_/X __dut__._1633_/X VGND VGND VPWR
+ VPWR __dut__._2874_/D sky130_fd_sc_hd__a21o_4
X__dut__._1565_ __dut__._1565_/A __dut__._2856_/Q VGND VGND VPWR VPWR __dut__._1565_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_58_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1496_ __dut__._1374_/Y mp[5] __dut__._1495_/X VGND VGND VPWR VPWR __dut__._1496_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2539__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1443__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1075__A __dut__.__uuf__._1640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3097_ __dut__._3102_/CLK __dut__._3097_/D __dut__._2521_/Y VGND VGND VPWR
+ VPWR __dut__._3097_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2117_ __dut__._2325_/A __dut__._2117_/B VGND VGND VPWR VPWR __dut__._2117_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2048_ __dut__._2412_/A1 prod[6] __dut__._2047_/X VGND VGND VPWR VPWR __dut__._3081_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_41_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2449__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_221_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1596__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2825__CLK __dut__._2846_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2352_ __dut__.__uuf__._2353_/CLK __dut__._2484_/X __dut__.__uuf__._1062_/X
+ VGND VGND VPWR VPWR prod[51] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1303_ __dut__.__uuf__._1300_/X __dut__.__uuf__._1302_/X __dut__._2353_/B
+ __dut__.__uuf__._1300_/X VGND VGND VPWR VPWR __dut__._2352_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._2283_ __dut__.__uuf__._2288_/CLK __dut__._2346_/X __dut__.__uuf__._1314_/X
+ VGND VGND VPWR VPWR __dut__._2347_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_99_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1234_ __dut__.__uuf__._1234_/A VGND VGND VPWR VPWR __dut__.__uuf__._1234_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_115_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1520__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1165_ __dut__.__uuf__._1175_/A VGND VGND VPWR VPWR __dut__.__uuf__._1165_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1096_ __dut__.__uuf__._1126_/A VGND VGND VPWR VPWR __dut__.__uuf__._1096_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2359__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._3020_ clkbuf_opt_2_tck/X __dut__._3020_/D __dut__._2598_/Y VGND VGND VPWR
+ VPWR __dut__._3020_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_91_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1998_ VGND VGND VPWR VPWR __dut__.__uuf__._1998_/HI tie[5] sky130_fd_sc_hd__conb_1
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_160_ _193_/B VGND VGND VPWR VPWR _172_/B sky130_fd_sc_hd__buf_2
XFILLER_155_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2804_ rst VGND VGND VPWR VPWR __dut__._2804_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2735_ rst VGND VGND VPWR VPWR __dut__._2735_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2666_ rst VGND VGND VPWR VPWR __dut__._2666_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1617_ __dut__._2105_/A __dut__._2869_/Q VGND VGND VPWR VPWR __dut__._1617_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2597_ rst VGND VGND VPWR VPWR __dut__._2597_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1548_ __dut__._1374_/Y mp[17] __dut__._1547_/X VGND VGND VPWR VPWR __dut__._1548_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_73_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1479_ __dut__._2509_/A __dut__._2836_/Q VGND VGND VPWR VPWR __dut__._1479_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_61_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1901__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2848__CLK __dut__._2860_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1533__A __dut__.__uuf__._1533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_289_ _290_/CLK _289_/D VGND VGND VPWR VPWR _289_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._2732__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0_tck_A clkbuf_3_1_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2451__B prod[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_171_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_269_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2179__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2058__A2 prod[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1921_ __dut__.__uuf__._1921_/A VGND VGND VPWR VPWR __dut__.__uuf__._1921_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1852_ __dut__._2187_/B __dut__._2193_/B VGND VGND VPWR VPWR __dut__.__uuf__._1853_/A
+ sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_4_11_0_tck_A clkbuf_3_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1783_ __dut__.__uuf__._1815_/A __dut__.__uuf__._1783_/B __dut__.__uuf__._1783_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1784_/A sky130_fd_sc_hd__or3_4
XFILLER_146_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2642__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2335_ __dut__.__uuf__._2364_/CLK __dut__._2450_/X __dut__.__uuf__._1113_/X
+ VGND VGND VPWR VPWR prod[34] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2520_ rst VGND VGND VPWR VPWR __dut__._2520_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2266_ __dut__.__uuf__._2291_/CLK __dut__._2312_/X __dut__.__uuf__._1402_/X
+ VGND VGND VPWR VPWR __dut__._2313_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1217_ __dut__._2373_/B VGND VGND VPWR VPWR __dut__.__uuf__._1248_/A
+ sky130_fd_sc_hd__inv_2
X__dut__._2451_ __dut__._2457_/A prod[34] VGND VGND VPWR VPWR __dut__._2451_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._2197_ __dut__.__uuf__._2230_/CLK __dut__._2174_/X __dut__.__uuf__._1606_/X
+ VGND VGND VPWR VPWR __dut__._2175_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1148_ __dut__.__uuf__._1147_/X __dut__.__uuf__._1144_/X prod[23]
+ prod[24] __dut__.__uuf__._1141_/X VGND VGND VPWR VPWR __dut__._2428_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1402_ __dut__._1418_/A1 __dut__._1400_/X __dut__._1401_/X VGND VGND VPWR
+ VPWR __dut__._2816_/D sky130_fd_sc_hd__a21o_4
XFILLER_142_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2382_ __dut__._2412_/A1 __dut__._2382_/A2 __dut__._2381_/X VGND VGND VPWR
+ VPWR __dut__._2382_/X sky130_fd_sc_hd__a21o_4
XFILLER_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1079_ __dut__.__uuf__._1087_/A VGND VGND VPWR VPWR __dut__.__uuf__._1079_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1721__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3003_ _306_/CLK __dut__._3003_/D __dut__._2615_/Y VGND VGND VPWR VPWR __dut__._3003_/Q
+ sky130_fd_sc_hd__dfrtp_4
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ _204_/Y _208_/X _211_/X _254_/Q _246_/Q VGND VGND VPWR VPWR tdo sky130_fd_sc_hd__a32o_4
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1980__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2552__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_143_ _295_/Q _296_/Q VGND VGND VPWR VPWR _220_/A sky130_fd_sc_hd__or2_4
XFILLER_109_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2718_ rst VGND VGND VPWR VPWR __dut__._2718_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2649_ rst VGND VGND VPWR VPWR __dut__._2649_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._1528__A __dut__.__uuf__._1549_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2727__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1631__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3026__CLK clkbuf_5_1_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1263__A __dut__.__uuf__._1533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2120_ VGND VGND VPWR VPWR __dut__.__uuf__._2120_/HI tie[127] sky130_fd_sc_hd__conb_1
XFILLER_130_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2051_ VGND VGND VPWR VPWR __dut__.__uuf__._2051_/HI tie[58] sky130_fd_sc_hd__conb_1
XFILLER_96_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2637__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1904_ __dut__.__uuf__._1904_/A VGND VGND VPWR VPWR __dut__.__uuf__._1952_/A
+ sky130_fd_sc_hd__buf_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1835_ __dut__.__uuf__._1835_/A VGND VGND VPWR VPWR __dut__.__uuf__._1837_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1766_ __dut__._2155_/B __dut__._2161_/B VGND VGND VPWR VPWR __dut__.__uuf__._1767_/A
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1962__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1951_ __dut__._2207_/A __dut__._3032_/Q VGND VGND VPWR VPWR __dut__._1951_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1697_ __dut__._1552_/X VGND VGND VPWR VPWR __dut__.__uuf__._1701_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1882_ __dut__._1882_/A1 tie[93] __dut__._1881_/X VGND VGND VPWR VPWR __dut__._2998_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2318_ __dut__.__uuf__._2328_/CLK __dut__._2416_/X __dut__.__uuf__._1165_/X
+ VGND VGND VPWR VPWR prod[17] sky130_fd_sc_hd__dfrtp_4
X__dut__._2503_ __dut__._2503_/A prod[60] VGND VGND VPWR VPWR __dut__._2503_/X sky130_fd_sc_hd__and2_4
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2249_ __dut__.__uuf__._2251_/CLK __dut__._2278_/X __dut__.__uuf__._1479_/X
+ VGND VGND VPWR VPWR __dut__._2279_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_153_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2434_ __dut__._2434_/A1 __dut__._2434_/A2 __dut__._2433_/X VGND VGND VPWR
+ VPWR __dut__._2434_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_72_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2365_ __dut__._2407_/A __dut__._2365_/B VGND VGND VPWR VPWR __dut__._2365_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._3049__CLK __dut__._3058_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2547__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2296_ __dut__._2296_/A1 __dut__._2296_/A2 __dut__._2295_/X VGND VGND VPWR
+ VPWR __dut__._2296_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1451__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2179__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_126_ _256_/D _258_/D VGND VGND VPWR VPWR _127_/D sky130_fd_sc_hd__and2_4
XFILLER_98_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_134_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1620_ __dut__.__uuf__._1621_/A VGND VGND VPWR VPWR __dut__.__uuf__._1620_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1944__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1551_ __dut__._1492_/X __dut__.__uuf__._1550_/X __dut__._2249_/B
+ __dut__.__uuf__._1534_/X VGND VGND VPWR VPWR __dut__.__uuf__._1551_/X sky130_fd_sc_hd__o22a_4
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1482_ __dut__.__uuf__._1463_/X __dut__.__uuf__._1480_/X __dut__._2279_/B
+ __dut__.__uuf__._1469_/X __dut__.__uuf__._1481_/X VGND VGND VPWR VPWR __dut__._2278_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2103_ VGND VGND VPWR VPWR __dut__.__uuf__._2103_/HI tie[110] sky130_fd_sc_hd__conb_1
XFILLER_131_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2034_ VGND VGND VPWR VPWR __dut__.__uuf__._2034_/HI tie[41] sky130_fd_sc_hd__conb_1
XFILLER_45_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2150_ __dut__._2208_/A1 __dut__._2150_/A2 __dut__._2149_/X VGND VGND VPWR
+ VPWR __dut__._2150_/X sky130_fd_sc_hd__a21o_4
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2367__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2081_ __dut__._2081_/A __dut__._3097_/Q VGND VGND VPWR VPWR __dut__._2081_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_80_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1818_ __dut__.__uuf__._1926_/A VGND VGND VPWR VPWR __dut__.__uuf__._1869_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_40_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1749_ __dut__.__uuf__._1704_/X __dut__.__uuf__._1747_/B __dut__.__uuf__._1747_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1750_/C sky130_fd_sc_hd__o21a_4
X__dut__._2983_ __dut__._2985_/CLK __dut__._2983_/D __dut__._2635_/Y VGND VGND VPWR
+ VPWR __dut__._2983_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1934_ __dut__._1942_/A1 tie[119] __dut__._1933_/X VGND VGND VPWR VPWR __dut__._3024_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1865_ __dut__._1881_/A __dut__._2989_/Q VGND VGND VPWR VPWR __dut__._1865_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2360__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1796_ __dut__._1830_/A1 tie[50] __dut__._1795_/X VGND VGND VPWR VPWR __dut__._2955_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_121_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_6_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2417_ __dut__._2417_/A prod[17] VGND VGND VPWR VPWR __dut__._2417_/X sky130_fd_sc_hd__and2_4
XFILLER_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2348_ __dut__._2368_/A1 __dut__._2348_/A2 __dut__._2347_/X VGND VGND VPWR
+ VPWR __dut__._2348_/X sky130_fd_sc_hd__a21o_4
XFILLER_73_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2279_ __dut__._2281_/A __dut__._2279_/B VGND VGND VPWR VPWR __dut__._2279_/X
+ sky130_fd_sc_hd__and2_4
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__282__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1210__A1 __dut__.__uuf__._1206_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2740__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_251_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1603_ __dut__.__uuf__._1603_/A VGND VGND VPWR VPWR __dut__.__uuf__._1628_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1534_ __dut__.__uuf__._1709_/A VGND VGND VPWR VPWR __dut__.__uuf__._1534_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2650__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1465_ __dut__.__uuf__._1550_/A VGND VGND VPWR VPWR __dut__.__uuf__._1465_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2342__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1650_ __dut__._2488_/A1 prod[42] __dut__._1649_/X VGND VGND VPWR VPWR __dut__._2882_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1396_ __dut__.__uuf__._1411_/A VGND VGND VPWR VPWR __dut__.__uuf__._1396_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1581_ __dut__._1589_/A __dut__._2860_/Q VGND VGND VPWR VPWR __dut__._1581_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2017_ VGND VGND VPWR VPWR __dut__.__uuf__._2017_/HI tie[24] sky130_fd_sc_hd__conb_1
XFILLER_85_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_6_0___dut__.__uuf__.__clk_source__ clkbuf_4_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2291_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_150_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2097__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2202_ __dut__._2202_/A1 __dut__._2202_/A2 __dut__._2201_/X VGND VGND VPWR
+ VPWR __dut__._2202_/X sky130_fd_sc_hd__a21o_4
X__dut__._2133_ __dut__._2141_/A __dut__._2133_/B VGND VGND VPWR VPWR __dut__._2133_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_35_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2881__CLK __dut__._3106_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2064_ __dut__._2412_/A1 prod[14] __dut__._2063_/X VGND VGND VPWR VPWR __dut__._3089_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1908__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1384__A2 mc[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2966_ __dut__._2985_/CLK __dut__._2966_/D __dut__._2652_/Y VGND VGND VPWR
+ VPWR __dut__._2966_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2560__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1917_ __dut__._2207_/A __dut__._3015_/Q VGND VGND VPWR VPWR __dut__._1917_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_141_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2897_ _306_/CLK __dut__._2897_/D __dut__._2721_/Y VGND VGND VPWR VPWR __dut__._2897_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_122_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1848_ __dut__._1848_/A1 tie[76] __dut__._1847_/X VGND VGND VPWR VPWR __dut__._2981_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_110_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1779_ __dut__._1779_/A __dut__._2946_/Q VGND VGND VPWR VPWR __dut__._1779_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2735__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_172 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1816_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_150 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2096_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_161 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1638_/A1 sky130_fd_sc_hd__buf_2
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_183 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._1382_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_194 psn_inst_psn_buff_201/A VGND VGND VPWR VPWR __dut__._1466_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_145_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_17 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2020_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_28 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1954_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_39 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2128_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_144_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2324__A1 __dut__._2332_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1250_ __dut__.__uuf__._1254_/A VGND VGND VPWR VPWR __dut__.__uuf__._1250_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1181_ __dut__.__uuf__._1177_/X __dut__.__uuf__._1173_/X prod[12]
+ prod[13] __dut__.__uuf__._1170_/X VGND VGND VPWR VPWR __dut__._2406_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_140_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_3_0_tck clkbuf_5_3_0_tck/A VGND VGND VPWR VPWR clkbuf_5_3_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2645__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2820_ __dut__._2509_/B __dut__._2820_/D __dut__._2798_/Y VGND VGND VPWR
+ VPWR __dut__._2820_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1517_ __dut__._1528_/X __dut__.__uuf__._1508_/X __dut__._2265_/B
+ __dut__.__uuf__._1513_/X VGND VGND VPWR VPWR __dut__.__uuf__._1517_/X sky130_fd_sc_hd__o22a_4
X__dut__._2751_ rst VGND VGND VPWR VPWR __dut__._2751_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1702_ __dut__._1714_/A1 tie[3] __dut__._1701_/X VGND VGND VPWR VPWR __dut__._2908_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2682_ rst VGND VGND VPWR VPWR __dut__._2682_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1448_ __dut__.__uuf__._1492_/A VGND VGND VPWR VPWR __dut__.__uuf__._1448_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1186__B1 prod[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1633_ __dut__._2197_/A __dut__._2873_/Q VGND VGND VPWR VPWR __dut__._1633_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1379_ __dut__._2325_/B VGND VGND VPWR VPWR __dut__.__uuf__._1379_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1564_ __dut__._1374_/Y mp[20] __dut__._1563_/X VGND VGND VPWR VPWR __dut__._1564_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1495_ __dut__._2509_/A __dut__._2840_/Q VGND VGND VPWR VPWR __dut__._1495_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2555__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3096_ __dut__._3096_/CLK __dut__._3096_/D __dut__._2522_/Y VGND VGND VPWR
+ VPWR __dut__._3096_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2116_ __dut__._2288_/A1 __dut__._2116_/A2 __dut__._2115_/X VGND VGND VPWR
+ VPWR __dut__._2116_/X sky130_fd_sc_hd__a21o_4
X__dut__._2047_ __dut__._2407_/A __dut__._3080_/Q VGND VGND VPWR VPWR __dut__._2047_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2949_ __dut__._2961_/CLK __dut__._2949_/D __dut__._2669_/Y VGND VGND VPWR
+ VPWR __dut__._2949_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2449__B prod[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2465__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_214_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1596__A2 mc[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2351_ __dut__.__uuf__._2353_/CLK __dut__._2482_/X __dut__.__uuf__._1064_/X
+ VGND VGND VPWR VPWR prod[50] sky130_fd_sc_hd__dfrtp_4
XFILLER_126_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1302_ __dut__.__uuf__._1301_/Y __dut__.__uuf__._1294_/X __dut__.__uuf__._1296_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1302_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._2282_ __dut__.__uuf__._2288_/CLK __dut__._2344_/X __dut__.__uuf__._1318_/X
+ VGND VGND VPWR VPWR __dut__._2345_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_114_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1233_ __dut__.__uuf__._1214_/A __dut__.__uuf__._1226_/X __dut__.__uuf__._1227_/X
+ __dut__._2381_/B __dut__.__uuf__._1232_/X VGND VGND VPWR VPWR __dut__._2380_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_115_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1183__A3 prod[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1520__A2 mp[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1164_ __dut__.__uuf__._1208_/A VGND VGND VPWR VPWR __dut__.__uuf__._1175_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_55_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1095_ __dut__.__uuf__._1101_/A VGND VGND VPWR VPWR __dut__.__uuf__._1095_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1176__A __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._3082__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1997_ VGND VGND VPWR VPWR __dut__.__uuf__._1997_/HI tie[4] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2375__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1904__A __dut__.__uuf__._1904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2803_ rst VGND VGND VPWR VPWR __dut__._2803_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1719__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2734_ rst VGND VGND VPWR VPWR __dut__._2734_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2665_ rst VGND VGND VPWR VPWR __dut__._2665_/Y sky130_fd_sc_hd__inv_2
X__dut__._2596_ rst VGND VGND VPWR VPWR __dut__._2596_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1616_ __dut__._1374_/Y start __dut__._1615_/X VGND VGND VPWR VPWR __dut__._1616_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_77_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1547_ __dut__._2509_/A __dut__._2853_/Q VGND VGND VPWR VPWR __dut__._1547_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1478_ __dut__._1478_/A1 __dut__._1476_/X __dut__._1477_/X VGND VGND VPWR
+ VPWR __dut__._2835_/D sky130_fd_sc_hd__a21o_4
XFILLER_61_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__311__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3079_ __dut__._3079_/CLK __dut__._3079_/D __dut__._2539_/Y VGND VGND VPWR
+ VPWR __dut__._3079_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_288_ _290_/CLK _288_/D VGND VGND VPWR VPWR _288_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_154_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_164_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1920_ __dut__.__uuf__._1920_/A VGND VGND VPWR VPWR __dut__.__uuf__._1923_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1851_ __dut__._1412_/X VGND VGND VPWR VPWR __dut__.__uuf__._1855_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1782_ __dut__.__uuf__._1759_/X __dut__.__uuf__._1780_/B __dut__.__uuf__._1780_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1783_/C sky130_fd_sc_hd__o21a_4
XFILLER_118_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1539__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2334_ __dut__.__uuf__._2334_/CLK __dut__._2448_/X __dut__.__uuf__._1117_/X
+ VGND VGND VPWR VPWR prod[33] sky130_fd_sc_hd__dfrtp_4
XFILLER_126_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2265_ __dut__.__uuf__._2291_/CLK __dut__._2310_/X __dut__.__uuf__._1407_/X
+ VGND VGND VPWR VPWR __dut__._2311_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_120_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1216_ __dut__.__uuf__._1234_/A VGND VGND VPWR VPWR __dut__.__uuf__._1216_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2450_ __dut__._2450_/A1 __dut__._2450_/A2 __dut__._2449_/X VGND VGND VPWR
+ VPWR __dut__._2450_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2196_ __dut__.__uuf__._2230_/CLK __dut__._2172_/X __dut__.__uuf__._1607_/X
+ VGND VGND VPWR VPWR __dut__._2173_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1401_ __dut__._2189_/A __dut__._2815_/Q VGND VGND VPWR VPWR __dut__._1401_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1147_ __dut__.__uuf__._1162_/A VGND VGND VPWR VPWR __dut__.__uuf__._1147_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2381_ __dut__._2407_/A __dut__._2381_/B VGND VGND VPWR VPWR __dut__._2381_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_142_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1078_ __dut__.__uuf__._1072_/X __dut__.__uuf__._1069_/X prod[47]
+ prod[48] __dut__.__uuf__._1066_/X VGND VGND VPWR VPWR __dut__._2476_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_83_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3002_ _306_/CLK __dut__._3002_/D __dut__._2616_/Y VGND VGND VPWR VPWR __dut__._3002_/Q
+ sky130_fd_sc_hd__dfrtp_4
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1634__A __dut__.__uuf__._1640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ _211_/A _211_/B VGND VGND VPWR VPWR _211_/X sky130_fd_sc_hd__or2_4
XFILLER_11_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_142_ _296_/Q VGND VGND VPWR VPWR _142_/Y sky130_fd_sc_hd__inv_2
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2717_ rst VGND VGND VPWR VPWR __dut__._2717_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2648_ rst VGND VGND VPWR VPWR __dut__._2648_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1496__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2579_ rst VGND VGND VPWR VPWR __dut__._2579_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1544__A __dut__.__uuf__._1563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1420__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2743__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_281_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2050_ VGND VGND VPWR VPWR __dut__.__uuf__._2050_/HI tie[57] sky130_fd_sc_hd__conb_1
XFILLER_57_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1903_ __dut__.__uuf__._1896_/A __dut__.__uuf__._1901_/B __dut__.__uuf__._1882_/X
+ VGND VGND VPWR VPWR __dut__._2202_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_80_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1834_ __dut__.__uuf__._1844_/A __dut__.__uuf__._1834_/B __dut__.__uuf__._1834_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1835_/A sky130_fd_sc_hd__or3_4
XANTENNA___dut__._2653__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1765_ __dut__._1380_/X VGND VGND VPWR VPWR __dut__.__uuf__._1769_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._1950_ __dut__._2172_/A1 tie[127] __dut__._1949_/X VGND VGND VPWR VPWR __dut__._3032_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1962__A2 tie[133] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1696_ __dut__.__uuf__._1689_/A __dut__.__uuf__._1694_/B __dut__.__uuf__._1661_/X
+ VGND VGND VPWR VPWR __dut__._2126_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1881_ __dut__._1881_/A __dut__._2997_/Q VGND VGND VPWR VPWR __dut__._1881_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_133_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2317_ __dut__.__uuf__._2328_/CLK __dut__._2414_/X __dut__.__uuf__._1167_/X
+ VGND VGND VPWR VPWR prod[16] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2838__CLK __dut__._2846_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2248_ __dut__.__uuf__._2251_/CLK __dut__._2276_/X __dut__.__uuf__._1485_/X
+ VGND VGND VPWR VPWR __dut__._2277_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2502_ __dut__._2502_/A1 __dut__._2502_/A2 __dut__._2501_/X VGND VGND VPWR
+ VPWR __dut__._2502_/X sky130_fd_sc_hd__a21o_4
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2179_ __dut__.__uuf__._2216_/CLK __dut__._2138_/X __dut__.__uuf__._1627_/X
+ VGND VGND VPWR VPWR __dut__._2139_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_48_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2433_ __dut__._2491_/A prod[25] VGND VGND VPWR VPWR __dut__._2433_/X sky130_fd_sc_hd__and2_4
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2364_ __dut__._2368_/A1 __dut__._2364_/A2 __dut__._2363_/X VGND VGND VPWR
+ VPWR __dut__._2364_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_65_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2295_ __dut__._2295_/A __dut__._2295_/B VGND VGND VPWR VPWR __dut__._2295_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1650__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2563__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1402__A1 __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_125_ _237_/A _138_/B VGND VGND VPWR VPWR _125_/X sky130_fd_sc_hd__and2_4
XFILLER_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1907__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2738__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2457__B prod[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_127_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2473__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1550_ __dut__.__uuf__._1550_/A VGND VGND VPWR VPWR __dut__.__uuf__._1550_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2273__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1481_ __dut__._1564_/X __dut__.__uuf__._1465_/X __dut__._2281_/B
+ __dut__.__uuf__._1470_/X VGND VGND VPWR VPWR __dut__.__uuf__._1481_/X sky130_fd_sc_hd__o22a_4
XFILLER_128_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2102_ VGND VGND VPWR VPWR __dut__.__uuf__._2102_/HI tie[109] sky130_fd_sc_hd__conb_1
XFILLER_131_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2033_ VGND VGND VPWR VPWR __dut__.__uuf__._2033_/HI tie[40] sky130_fd_sc_hd__conb_1
XFILLER_29_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2648__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2080_ __dut__._2428_/A1 prod[22] __dut__._2079_/X VGND VGND VPWR VPWR __dut__._3097_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1632__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1817_ __dut__.__uuf__._1809_/A __dut__.__uuf__._1815_/B __dut__.__uuf__._1774_/X
+ VGND VGND VPWR VPWR __dut__._2170_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_138_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1748_ __dut__.__uuf__._1748_/A VGND VGND VPWR VPWR __dut__.__uuf__._1750_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._2982_ __dut__._2985_/CLK __dut__._2982_/D __dut__._2636_/Y VGND VGND VPWR
+ VPWR __dut__._2982_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1933_ __dut__._2207_/A __dut__._3023_/Q VGND VGND VPWR VPWR __dut__._1933_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1679_ __dut__._2123_/B __dut__._2129_/B __dut__.__uuf__._1678_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1680_/C sky130_fd_sc_hd__o21ai_4
XFILLER_153_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1864_ __dut__._1864_/A1 tie[84] __dut__._1863_/X VGND VGND VPWR VPWR __dut__._2989_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1727__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3016__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1795_ __dut__._1797_/A __dut__._2954_/Q VGND VGND VPWR VPWR __dut__._1795_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2416_ __dut__._2422_/A1 __dut__._2416_/A2 __dut__._2415_/X VGND VGND VPWR
+ VPWR __dut__._2416_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2558__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2347_ __dut__._2407_/A __dut__._2347_/B VGND VGND VPWR VPWR __dut__._2347_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2278_ __dut__._2278_/A1 __dut__._2278_/A2 __dut__._2277_/X VGND VGND VPWR
+ VPWR __dut__._2278_/X sky130_fd_sc_hd__a21o_4
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._2296__CLK __dut__.__uuf__._2303_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1637__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_244_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1372__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1602_ __dut__.__uuf__._1602_/A VGND VGND VPWR VPWR __dut__.__uuf__._1602_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1378__B1 __dut__._1377_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1533_ __dut__.__uuf__._1533_/A VGND VGND VPWR VPWR __dut__.__uuf__._1533_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1464_ __dut__.__uuf__._1464_/A VGND VGND VPWR VPWR __dut__.__uuf__._1550_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_104_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1547__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1395_ __dut__.__uuf__._1389_/X __dut__.__uuf__._1394_/X __dut__._2317_/B
+ __dut__.__uuf__._1389_/X VGND VGND VPWR VPWR __dut__._2316_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1580_ __dut__._1374_/Y mp[24] __dut__._1579_/X VGND VGND VPWR VPWR __dut__._1580_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_69_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2169__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2016_ VGND VGND VPWR VPWR __dut__.__uuf__._2016_/HI tie[23] sky130_fd_sc_hd__conb_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2201_ __dut__._2207_/A __dut__._2201_/B VGND VGND VPWR VPWR __dut__._2201_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_27_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2132_ __dut__._2132_/A1 __dut__._2132_/A2 __dut__._2131_/X VGND VGND VPWR
+ VPWR __dut__._2132_/X sky130_fd_sc_hd__a21o_4
X__dut__._2063_ __dut__._2407_/A __dut__._3088_/Q VGND VGND VPWR VPWR __dut__._2063_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_28_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2965_ __dut__._2985_/CLK __dut__._2965_/D __dut__._2653_/Y VGND VGND VPWR
+ VPWR __dut__._2965_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1916_ __dut__._1916_/A1 tie[110] __dut__._1915_/X VGND VGND VPWR VPWR __dut__._3015_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2896_ _306_/CLK __dut__._2896_/D __dut__._2722_/Y VGND VGND VPWR VPWR __dut__._2896_/Q
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1457__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1847_ __dut__._1881_/A __dut__._2980_/Q VGND VGND VPWR VPWR __dut__._1847_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1778_ __dut__._1780_/A1 tie[41] __dut__._1777_/X VGND VGND VPWR VPWR __dut__._2946_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_140 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2430_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_173 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2376_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_151 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2444_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_162 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2506_/A1 sky130_fd_sc_hd__buf_2
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_184 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._1698_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_195 psn_inst_psn_buff_201/A VGND VGND VPWR VPWR __dut__._2212_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_18 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2018_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_29 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1952_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2751__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1180_ __dut__.__uuf__._1191_/A VGND VGND VPWR VPWR __dut__.__uuf__._1180_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_140_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2088__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1516_ __dut__.__uuf__._1522_/A VGND VGND VPWR VPWR __dut__.__uuf__._1516_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2661__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2750_ rst VGND VGND VPWR VPWR __dut__._2750_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1701_ __dut__._2189_/A __dut__._2907_/Q VGND VGND VPWR VPWR __dut__._1701_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2681_ rst VGND VGND VPWR VPWR __dut__._2681_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1447_ __dut__.__uuf__._1447_/A VGND VGND VPWR VPWR __dut__.__uuf__._1447_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_145_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1378_ __dut__.__uuf__._1378_/A VGND VGND VPWR VPWR __dut__.__uuf__._1378_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1632_ __dut__._1374_/Y mc[9] __dut__._1631_/X VGND VGND VPWR VPWR __dut__._1632_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_77_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__272__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1563_ __dut__._2509_/A __dut__._2857_/Q VGND VGND VPWR VPWR __dut__._1563_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1494_ __dut__._2262_/A1 __dut__._1492_/X __dut__._1493_/X VGND VGND VPWR
+ VPWR __dut__._2839_/D sky130_fd_sc_hd__a21o_4
XFILLER_73_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2115_ __dut__._2325_/A __dut__._2115_/B VGND VGND VPWR VPWR __dut__._2115_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._3095_ __dut__._3096_/CLK __dut__._3095_/D __dut__._2523_/Y VGND VGND VPWR
+ VPWR __dut__._3095_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2046_ __dut__._2412_/A1 prod[5] __dut__._2045_/X VGND VGND VPWR VPWR __dut__._3080_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_110_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2571__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2948_ __dut__._2961_/CLK __dut__._2948_/D __dut__._2670_/Y VGND VGND VPWR
+ VPWR __dut__._2948_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2879_ __dut__._3106_/CLK __dut__._2879_/D __dut__._2739_/Y VGND VGND VPWR
+ VPWR __dut__._2879_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1915__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_19_0_tck clkbuf_4_9_0_tck/X VGND VGND VPWR VPWR __dut__._3093_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2490__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2746__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_207_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2481__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2350_ __dut__.__uuf__._2353_/CLK __dut__._2480_/X __dut__.__uuf__._1068_/X
+ VGND VGND VPWR VPWR prod[49] sky130_fd_sc_hd__dfrtp_4
XFILLER_132_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2281_ __dut__.__uuf__._2288_/CLK __dut__._2342_/X __dut__.__uuf__._1325_/X
+ VGND VGND VPWR VPWR __dut__._2343_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1301_ __dut__._2355_/B VGND VGND VPWR VPWR __dut__.__uuf__._1301_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_113_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1232_ __dut__.__uuf__._1414_/A VGND VGND VPWR VPWR __dut__.__uuf__._1232_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_141_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1163_ __dut__.__uuf__._1162_/X __dut__.__uuf__._1159_/X prod[18]
+ prod[19] __dut__.__uuf__._1156_/X VGND VGND VPWR VPWR __dut__._2418_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._2871__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1094_ __dut__.__uuf__._1088_/X __dut__.__uuf__._1085_/X prod[41]
+ prod[42] __dut__.__uuf__._1082_/X VGND VGND VPWR VPWR __dut__._2464_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_95_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2207__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2656__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1996_ VGND VGND VPWR VPWR __dut__.__uuf__._1996_/HI tie[3] sky130_fd_sc_hd__conb_1
XANTENNA___dut__.__uuf__._1192__A __dut__.__uuf__._1463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2802_ rst VGND VGND VPWR VPWR __dut__._2802_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2733_ rst VGND VGND VPWR VPWR __dut__._2733_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1735__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2664_ rst VGND VGND VPWR VPWR __dut__._2664_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2595_ rst VGND VGND VPWR VPWR __dut__._2595_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_95_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1615_ __dut__._2509_/A __dut__._2870_/Q VGND VGND VPWR VPWR __dut__._1615_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1546_ __dut__._1562_/A1 __dut__._1544_/X __dut__._1545_/X VGND VGND VPWR
+ VPWR __dut__._2852_/D sky130_fd_sc_hd__a21o_4
XFILLER_92_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2472__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1477_ __dut__._2281_/A __dut__._2834_/Q VGND VGND VPWR VPWR __dut__._1477_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2566__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3078_ __dut__._3093_/CLK __dut__._3078_/D __dut__._2540_/Y VGND VGND VPWR
+ VPWR __dut__._3078_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2029_ __dut__._2207_/A __dut__._3071_/Q VGND VGND VPWR VPWR __dut__._2029_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_81_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_287_ _290_/CLK _287_/D VGND VGND VPWR VPWR _287_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_154_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2894__CLK __dut__._3106_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_2_0_tck clkbuf_5_3_0_tck/A VGND VGND VPWR VPWR clkbuf_5_2_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1645__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_157_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1850_ __dut__.__uuf__._1904_/A VGND VGND VPWR VPWR __dut__.__uuf__._1898_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1781_ __dut__.__uuf__._1781_/A VGND VGND VPWR VPWR __dut__.__uuf__._1783_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_137_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2333_ __dut__.__uuf__._2334_/CLK __dut__._2446_/X __dut__.__uuf__._1121_/X
+ VGND VGND VPWR VPWR prod[32] sky130_fd_sc_hd__dfrtp_4
XFILLER_102_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2264_ __dut__.__uuf__._2291_/CLK __dut__._2308_/X __dut__.__uuf__._1411_/X
+ VGND VGND VPWR VPWR __dut__._2309_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_113_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1555__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1215_ __dut__.__uuf__._1206_/X __dut__.__uuf__._1203_/X prod[0]
+ prod[1] __dut__.__uuf__._1214_/X VGND VGND VPWR VPWR __dut__._2382_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._2195_ __dut__.__uuf__._2230_/CLK __dut__._2170_/X __dut__.__uuf__._1608_/X
+ VGND VGND VPWR VPWR __dut__._2171_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1146_ __dut__.__uuf__._1146_/A VGND VGND VPWR VPWR __dut__.__uuf__._1146_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1400_ __dut__._1374_/Y mc[15] __dut__._1399_/X VGND VGND VPWR VPWR __dut__._1400_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2380_ __dut__._2412_/A1 __dut__._2380_/A2 __dut__._2379_/X VGND VGND VPWR
+ VPWR __dut__._2380_/X sky130_fd_sc_hd__a21o_4
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1077_ __dut__.__uuf__._1087_/A VGND VGND VPWR VPWR __dut__.__uuf__._1077_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3001_ __dut__._3102_/CLK __dut__._3001_/D __dut__._2617_/Y VGND VGND VPWR
+ VPWR __dut__._3001_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_210_ _209_/Y _210_/A2 _247_/Q _253_/Q VGND VGND VPWR VPWR _211_/B sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1979_ __dut__._2235_/B __dut__._2117_/B VGND VGND VPWR VPWR __dut__.__uuf__._1980_/A
+ sky130_fd_sc_hd__and2_4
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_141_ _295_/Q VGND VGND VPWR VPWR _239_/A sky130_fd_sc_hd__buf_2
XFILLER_137_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_psn_inst_psn_buff_10_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2716_ rst VGND VGND VPWR VPWR __dut__._2716_/Y sky130_fd_sc_hd__inv_2
X__dut__._2647_ rst VGND VGND VPWR VPWR __dut__._2647_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1465__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1496__A2 mp[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2578_ rst VGND VGND VPWR VPWR __dut__._2578_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1529_ __dut__._1557_/A __dut__._2847_/Q VGND VGND VPWR VPWR __dut__._1529_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_19_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1420__A2 mc[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3072__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_274_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1902_ __dut__.__uuf__._1902_/A VGND VGND VPWR VPWR __dut__._2204_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_80_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1833_ __dut__._2179_/B __dut__._2185_/B __dut__.__uuf__._1832_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1834_/C sky130_fd_sc_hd__o21ai_4
XFILLER_40_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1764_ __dut__.__uuf__._1926_/A VGND VGND VPWR VPWR __dut__.__uuf__._1815_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_119_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1695_ __dut__.__uuf__._1695_/A VGND VGND VPWR VPWR __dut__._2128_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_118_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_9_0_tck clkbuf_4_9_0_tck/A VGND VGND VPWR VPWR clkbuf_4_9_0_tck/X sky130_fd_sc_hd__clkbuf_1
X__dut__._1880_ __dut__._1880_/A1 tie[92] __dut__._1879_/X VGND VGND VPWR VPWR __dut__._2997_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2316_ __dut__.__uuf__._2358_/CLK __dut__._2412_/X __dut__.__uuf__._1169_/X
+ VGND VGND VPWR VPWR prod[15] sky130_fd_sc_hd__dfrtp_4
XFILLER_121_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2247_ __dut__.__uuf__._2251_/CLK __dut__._2274_/X __dut__.__uuf__._1490_/X
+ VGND VGND VPWR VPWR __dut__._2275_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2501_ __dut__._2501_/A prod[59] VGND VGND VPWR VPWR __dut__._2501_/X sky130_fd_sc_hd__and2_4
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2178_ __dut__.__uuf__._2225_/CLK __dut__._2136_/X __dut__.__uuf__._1629_/X
+ VGND VGND VPWR VPWR __dut__._2137_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2432_ __dut__._2432_/A1 __dut__._2432_/A2 __dut__._2431_/X VGND VGND VPWR
+ VPWR __dut__._2432_/X sky130_fd_sc_hd__a21o_4
XFILLER_101_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1129_ __dut__.__uuf__._1173_/A VGND VGND VPWR VPWR __dut__.__uuf__._1129_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2363_ __dut__._2407_/A __dut__._2363_/B VGND VGND VPWR VPWR __dut__._2363_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_90_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2294_ __dut__._2294_/A1 __dut__._2294_/A2 __dut__._2293_/X VGND VGND VPWR
+ VPWR __dut__._2294_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_58_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1402__A2 __dut__._1400_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_124_ _291_/Q VGND VGND VPWR VPWR _138_/B sky130_fd_sc_hd__inv_2
XFILLER_152_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1923__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2754__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1480_ __dut__.__uuf__._1480_/A VGND VGND VPWR VPWR __dut__.__uuf__._1480_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2101_ VGND VGND VPWR VPWR __dut__.__uuf__._2101_/HI tie[108] sky130_fd_sc_hd__conb_1
XFILLER_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2032_ VGND VGND VPWR VPWR __dut__.__uuf__._2032_/HI tie[39] sky130_fd_sc_hd__conb_1
XFILLER_97_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1833__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1632__A2 mc[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2664__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1816_ __dut__.__uuf__._1816_/A VGND VGND VPWR VPWR __dut__._2172_/A2
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._1047__A3 prod[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1396__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1747_ __dut__.__uuf__._1790_/A __dut__.__uuf__._1747_/B __dut__.__uuf__._1747_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1748_/A sky130_fd_sc_hd__or3_4
X__dut__._2981_ __dut__._2985_/CLK __dut__._2981_/D __dut__._2637_/Y VGND VGND VPWR
+ VPWR __dut__._2981_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1932_ __dut__._1932_/A1 tie[118] __dut__._1931_/X VGND VGND VPWR VPWR __dut__._3023_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_153_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1678_ __dut__.__uuf__._1678_/A VGND VGND VPWR VPWR __dut__.__uuf__._1678_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_134_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1863_ __dut__._1881_/A __dut__._2988_/Q VGND VGND VPWR VPWR __dut__._1863_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1794_ __dut__._1830_/A1 tie[49] __dut__._1793_/X VGND VGND VPWR VPWR __dut__._2954_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_121_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2415_ __dut__._2415_/A prod[16] VGND VGND VPWR VPWR __dut__._2415_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1743__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2346_ __dut__._2368_/A1 __dut__._2346_/A2 __dut__._2345_/X VGND VGND VPWR
+ VPWR __dut__._2346_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2277_ __dut__._2281_/A __dut__._2277_/B VGND VGND VPWR VPWR __dut__._2277_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2574__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2749__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1653__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_237_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__.__uuf__._2240__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2828__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1601_ __dut__.__uuf__._1602_/A VGND VGND VPWR VPWR __dut__.__uuf__._1601_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_148_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1532_ __dut__.__uuf__._1543_/A VGND VGND VPWR VPWR __dut__.__uuf__._1532_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_116_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1463_ __dut__.__uuf__._1463_/A VGND VGND VPWR VPWR __dut__.__uuf__._1463_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_104_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1394_ __dut__.__uuf__._1393_/Y __dut__.__uuf__._1373_/X __dut__.__uuf__._1374_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1394_/X sky130_fd_sc_hd__o21a_4
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2659__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2015_ VGND VGND VPWR VPWR __dut__.__uuf__._2015_/HI tie[22] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._1563__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2200_ __dut__._2200_/A1 __dut__._2200_/A2 __dut__._2199_/X VGND VGND VPWR
+ VPWR __dut__._2200_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2131_ __dut__._2141_/A __dut__._2131_/B VGND VGND VPWR VPWR __dut__._2131_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_53_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2062_ __dut__._2412_/A1 prod[13] __dut__._2061_/X VGND VGND VPWR VPWR __dut__._3088_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_43_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2964_ __dut__._2985_/CLK __dut__._2964_/D __dut__._2654_/Y VGND VGND VPWR
+ VPWR __dut__._2964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1915_ __dut__._2005_/A __dut__._3014_/Q VGND VGND VPWR VPWR __dut__._1915_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2895_ __dut__._3106_/CLK __dut__._2895_/D __dut__._2723_/Y VGND VGND VPWR
+ VPWR __dut__._2895_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1846_ __dut__._1846_/A1 tie[75] __dut__._1845_/X VGND VGND VPWR VPWR __dut__._2980_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1777_ __dut__._1777_/A __dut__._2945_/Q VGND VGND VPWR VPWR __dut__._1777_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2569__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__305__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2329_ __dut__._2407_/A __dut__._2329_/B VGND VGND VPWR VPWR __dut__._2329_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_90_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1664__B1 __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_130 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1880_/A1 sky130_fd_sc_hd__buf_2
XFILLER_32_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_141 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2432_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_152 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2446_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_163 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2508_/A1 sky130_fd_sc_hd__buf_2
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_185 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._1696_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_174 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2278_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_196 psn_inst_psn_buff_201/A VGND VGND VPWR VPWR __dut__._2204_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_19 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._2016_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_145_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1532__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2479__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1383__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1515_ __dut__.__uuf__._1507_/X __dut__.__uuf__._1502_/X __dut__._2265_/B
+ __dut__.__uuf__._1512_/X __dut__.__uuf__._1514_/X VGND VGND VPWR VPWR __dut__._2264_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_135_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1700_ __dut__._1714_/A1 tie[2] __dut__._1699_/X VGND VGND VPWR VPWR __dut__._2907_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2680_ rst VGND VGND VPWR VPWR __dut__._2680_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1446_ __dut__.__uuf__._1446_/A VGND VGND VPWR VPWR __dut__.__uuf__._1447_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_145_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1377_ __dut__.__uuf__._1386_/A VGND VGND VPWR VPWR __dut__.__uuf__._1377_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1631_ __dut__._2509_/A __dut__._2874_/Q VGND VGND VPWR VPWR __dut__._1631_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1562_ __dut__._1562_/A1 __dut__._1560_/X __dut__._1561_/X VGND VGND VPWR
+ VPWR __dut__._2856_/D sky130_fd_sc_hd__a21o_4
XFILLER_100_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1493_ __dut__._1493_/A __dut__._2838_/Q VGND VGND VPWR VPWR __dut__._1493_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2114_ __dut__._2288_/A1 __dut__._2114_/A2 __dut__._2113_/X VGND VGND VPWR
+ VPWR __dut__._2114_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_40_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._3094_ __dut__._3096_/CLK __dut__._3094_/D __dut__._2524_/Y VGND VGND VPWR
+ VPWR __dut__._3094_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2045_ __dut__._2407_/A __dut__._3079_/Q VGND VGND VPWR VPWR __dut__._2045_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2947_ __dut__._2961_/CLK __dut__._2947_/D __dut__._2671_/Y VGND VGND VPWR
+ VPWR __dut__._2947_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_142_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2878_ __dut__._3109_/CLK __dut__._2878_/D __dut__._2740_/Y VGND VGND VPWR
+ VPWR __dut__._2878_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1829_ __dut__._1829_/A __dut__._2971_/Q VGND VGND VPWR VPWR __dut__._1829_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_96_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1828__A __dut__.__uuf__._1828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1931__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1563__A __dut__.__uuf__._1563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3029__CLK clkbuf_5_1_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2762__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_102_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__298__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2280_ __dut__.__uuf__._2288_/CLK __dut__._2340_/X __dut__.__uuf__._1331_/X
+ VGND VGND VPWR VPWR __dut__._2341_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1300_ __dut__.__uuf__._1311_/A VGND VGND VPWR VPWR __dut__.__uuf__._1300_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1231_ __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR __dut__.__uuf__._1414_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_141_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1162_ __dut__.__uuf__._1162_/A VGND VGND VPWR VPWR __dut__.__uuf__._1162_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1093_ __dut__.__uuf__._1101_/A VGND VGND VPWR VPWR __dut__.__uuf__._1093_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1841__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1995_ VGND VGND VPWR VPWR __dut__.__uuf__._1995_/HI tie[2] sky130_fd_sc_hd__conb_1
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1992__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2672__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2801_ rst VGND VGND VPWR VPWR __dut__._2801_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2732_ rst VGND VGND VPWR VPWR __dut__._2732_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1429_ __dut__.__uuf__._1255_/X __dut__.__uuf__._1428_/X __dut__._2303_/B
+ __dut__.__uuf__._1255_/X VGND VGND VPWR VPWR __dut__._2302_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_78_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2663_ rst VGND VGND VPWR VPWR __dut__._2663_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1614_ __dut__._2376_/A1 __dut__._1612_/X __dut__._1613_/X VGND VGND VPWR
+ VPWR __dut__._2869_/D sky130_fd_sc_hd__a21o_4
X__dut__._2594_ rst VGND VGND VPWR VPWR __dut__._2594_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_88_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1545_ __dut__._1557_/A __dut__._2851_/Q VGND VGND VPWR VPWR __dut__._1545_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1751__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1476_ __dut__._1374_/Y mp[0] __dut__._1475_/X VGND VGND VPWR VPWR __dut__._1476_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_73_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3077_ __dut__._3079_/CLK __dut__._3077_/D __dut__._2541_/Y VGND VGND VPWR
+ VPWR __dut__._3077_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._2301__CLK __dut__.__uuf__._2303_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2028_ __dut__._2028_/A1 tie[166] __dut__._2027_/X VGND VGND VPWR VPWR __dut__._3071_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2582__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_286_ _290_/CLK _286_/D VGND VGND VPWR VPWR _286_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_154_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2160__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1661__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2757__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1293__A __dut__.__uuf__._1709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1780_ __dut__.__uuf__._1790_/A __dut__.__uuf__._1780_/B __dut__.__uuf__._1780_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1781_/A sky130_fd_sc_hd__or3_4
XANTENNA___dut__._1974__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2332_ __dut__.__uuf__._2358_/CLK __dut__._2444_/X __dut__.__uuf__._1123_/X
+ VGND VGND VPWR VPWR prod[31] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2263_ __dut__.__uuf__._2293_/CLK __dut__._2306_/X __dut__.__uuf__._1417_/X
+ VGND VGND VPWR VPWR __dut__._2307_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_87_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1214_ __dut__.__uuf__._1214_/A VGND VGND VPWR VPWR __dut__.__uuf__._1214_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2194_ __dut__.__uuf__._2230_/CLK __dut__._2168_/X __dut__.__uuf__._1609_/X
+ VGND VGND VPWR VPWR __dut__._2169_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_75_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1145_ __dut__.__uuf__._1132_/X __dut__.__uuf__._1144_/X prod[24]
+ prod[25] __dut__.__uuf__._1141_/X VGND VGND VPWR VPWR __dut__._2430_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1076_ __dut__.__uuf__._1134_/A VGND VGND VPWR VPWR __dut__.__uuf__._1087_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1571__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2667__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3000_ __dut__._3096_/CLK __dut__._3000_/D __dut__._2618_/Y VGND VGND VPWR
+ VPWR __dut__._3000_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1978_ __dut__._1468_/X VGND VGND VPWR VPWR __dut__.__uuf__._1982_/B
+ sky130_fd_sc_hd__inv_2
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_140_ _140_/A VGND VGND VPWR VPWR _311_/D sky130_fd_sc_hd__inv_2
Xclkbuf_5_18_0_tck clkbuf_4_9_0_tck/X VGND VGND VPWR VPWR __dut__._3096_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2390__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2715_ rst VGND VGND VPWR VPWR __dut__._2715_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2646_ rst VGND VGND VPWR VPWR __dut__._2646_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2577_ rst VGND VGND VPWR VPWR __dut__._2577_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2577__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1528_ __dut__._1374_/Y mp[12] __dut__._1527_/X VGND VGND VPWR VPWR __dut__._1528_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1459_ __dut__._2509_/A __dut__._2831_/Q VGND VGND VPWR VPWR __dut__._1459_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_34_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__285__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_269_ _274_/CLK _269_/D VGND VGND VPWR VPWR _269_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_267_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1375__B __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1391__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2487__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1901_ __dut__.__uuf__._1923_/A __dut__.__uuf__._1901_/B __dut__.__uuf__._1901_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1902_/A sky130_fd_sc_hd__or3_4
XFILLER_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1832_ __dut__.__uuf__._1832_/A VGND VGND VPWR VPWR __dut__.__uuf__._1832_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_80_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1763_ __dut__.__uuf__._1755_/A __dut__.__uuf__._1761_/B __dut__.__uuf__._1720_/X
+ VGND VGND VPWR VPWR __dut__._2150_/A2 sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1694_ __dut__.__uuf__._1706_/A __dut__.__uuf__._1694_/B __dut__.__uuf__._1694_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1695_/A sky130_fd_sc_hd__or3_4
XFILLER_133_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2315_ __dut__.__uuf__._2358_/CLK __dut__._2410_/X __dut__.__uuf__._1172_/X
+ VGND VGND VPWR VPWR prod[14] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2124__A1 __dut__._2332_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2246_ __dut__.__uuf__._2251_/CLK __dut__._2272_/X __dut__.__uuf__._1495_/X
+ VGND VGND VPWR VPWR __dut__._2273_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2500_ __dut__._2502_/A1 __dut__._2500_/A2 __dut__._2499_/X VGND VGND VPWR
+ VPWR __dut__._2500_/X sky130_fd_sc_hd__a21o_4
XFILLER_102_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2431_ __dut__._2431_/A prod[24] VGND VGND VPWR VPWR __dut__._2431_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._2177_ __dut__.__uuf__._2225_/CLK __dut__._2134_/X __dut__.__uuf__._1630_/X
+ VGND VGND VPWR VPWR __dut__._2135_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1128_ __dut__.__uuf__._1131_/A VGND VGND VPWR VPWR __dut__.__uuf__._1128_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2397__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2362_ __dut__._2368_/A1 __dut__._2362_/A2 __dut__._2361_/X VGND VGND VPWR
+ VPWR __dut__._2362_/X sky130_fd_sc_hd__a21o_4
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2293_ __dut__._2293_/A __dut__._2293_/B VGND VGND VPWR VPWR __dut__._2293_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1059_ __dut__.__uuf__._1992_/A VGND VGND VPWR VPWR __dut__.__uuf__._1071_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_71_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2884__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_1_0_tck clkbuf_5_1_0_tck/A VGND VGND VPWR VPWR clkbuf_5_1_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__.__uuf__._1661__A __dut__.__uuf__._1828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_123_ _314_/Q VGND VGND VPWR VPWR _237_/A sky130_fd_sc_hd__inv_2
XFILLER_137_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2629_ rst VGND VGND VPWR VPWR __dut__._2629_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0___dut__.__uuf__.__clk_source__ clkbuf_2_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2770__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2354__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2100_ VGND VGND VPWR VPWR __dut__.__uuf__._2100_/HI tie[107] sky130_fd_sc_hd__conb_1
XFILLER_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2031_ VGND VGND VPWR VPWR __dut__.__uuf__._2031_/HI tie[38] sky130_fd_sc_hd__conb_1
XFILLER_97_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1815_ __dut__.__uuf__._1815_/A __dut__.__uuf__._1815_/B __dut__.__uuf__._1815_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1816_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1746_ __dut__._2147_/B __dut__._2153_/B __dut__.__uuf__._1745_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1747_/C sky130_fd_sc_hd__o21ai_4
XANTENNA___dut__._1396__A2 mc[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2980_ __dut__._3079_/CLK __dut__._2980_/D __dut__._2638_/Y VGND VGND VPWR
+ VPWR __dut__._2980_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1931_ __dut__._2207_/A __dut__._3022_/Q VGND VGND VPWR VPWR __dut__._1931_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_153_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1677_ __dut__._2123_/B __dut__._2129_/B VGND VGND VPWR VPWR __dut__.__uuf__._1678_/A
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2680__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1862_ __dut__._1864_/A1 tie[83] __dut__._1861_/X VGND VGND VPWR VPWR __dut__._2988_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1793_ __dut__._1797_/A __dut__._2953_/Q VGND VGND VPWR VPWR __dut__._1793_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2229_ __dut__.__uuf__._2230_/CLK __dut__._2238_/X __dut__.__uuf__._1562_/X
+ VGND VGND VPWR VPWR __dut__._2239_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2414_ __dut__._2422_/A1 __dut__._2414_/A2 __dut__._2413_/X VGND VGND VPWR
+ VPWR __dut__._2414_/X sky130_fd_sc_hd__a21o_4
XFILLER_91_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_70_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2345_ __dut__._2407_/A __dut__._2345_/B VGND VGND VPWR VPWR __dut__._2345_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2276_ __dut__._2278_/A1 __dut__._2276_/A2 __dut__._2275_/X VGND VGND VPWR
+ VPWR __dut__._2276_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._3062__CLK clkbuf_5_6_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2590__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2192__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2336__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0_tck clkbuf_4_9_0_tck/A VGND VGND VPWR VPWR clkbuf_4_8_0_tck/X sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._2765__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_132_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1682__A1 __dut__.__uuf__._1261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1600_ __dut__.__uuf__._1602_/A VGND VGND VPWR VPWR __dut__.__uuf__._1600_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1531_ __dut__.__uuf__._1528_/X __dut__.__uuf__._1523_/X __dut__._2257_/B
+ __dut__.__uuf__._1512_/X __dut__.__uuf__._1530_/X VGND VGND VPWR VPWR __dut__._2256_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_144_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1198__B1 prod[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1462_ __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR __dut__.__uuf__._1462_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2005__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1393_ __dut__._2319_/B VGND VGND VPWR VPWR __dut__.__uuf__._1393_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2014_ VGND VGND VPWR VPWR __dut__.__uuf__._2014_/HI tie[21] sky130_fd_sc_hd__conb_1
XFILLER_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._3085__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2130_ __dut__._2130_/A1 __dut__._2130_/A2 __dut__._2129_/X VGND VGND VPWR
+ VPWR __dut__._2130_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2675__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1122__B1 prod[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2061_ __dut__._2407_/A __dut__._3087_/Q VGND VGND VPWR VPWR __dut__._2061_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1729_ __dut__.__uuf__._1761_/A __dut__.__uuf__._1729_/B __dut__.__uuf__._1729_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1730_/A sky130_fd_sc_hd__or3_4
X__dut__._2963_ __dut__._3079_/CLK __dut__._2963_/D __dut__._2655_/Y VGND VGND VPWR
+ VPWR __dut__._2963_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1914_ __dut__._2004_/A1 tie[109] __dut__._1913_/X VGND VGND VPWR VPWR __dut__._3014_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2894_ __dut__._3106_/CLK __dut__._2894_/D __dut__._2724_/Y VGND VGND VPWR
+ VPWR __dut__._2894_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1845_ __dut__._1881_/A __dut__._2979_/Q VGND VGND VPWR VPWR __dut__._1845_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1776_ __dut__._1780_/A1 tie[40] __dut__._1775_/X VGND VGND VPWR VPWR __dut__._2945_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_4_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2328_ __dut__._2332_/A1 __dut__._2328_/A2 __dut__._2327_/X VGND VGND VPWR
+ VPWR __dut__._2328_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2585__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2259_ __dut__._2259_/A __dut__._2259_/B VGND VGND VPWR VPWR __dut__._2259_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_120 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1846_/A1 sky130_fd_sc_hd__buf_2
XFILLER_32_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2006__B1 __dut__._2005_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_142 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2488_/A1 sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_131 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1882_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_153 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2452_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_164 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1690_/A1 sky130_fd_sc_hd__buf_2
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_186 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._1726_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_175 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1490_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_197 psn_inst_psn_buff_201/A VGND VGND VPWR VPWR __dut__._2202_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1929__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1532__A2 mp[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1839__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1514_ __dut__._1532_/X __dut__.__uuf__._1508_/X __dut__._2267_/B
+ __dut__.__uuf__._1513_/X VGND VGND VPWR VPWR __dut__.__uuf__._1514_/X sky130_fd_sc_hd__o22a_4
XFILLER_135_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1445_ __dut__.__uuf__._1457_/A VGND VGND VPWR VPWR __dut__.__uuf__._1445_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1186__A3 prod[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1376_ __dut__.__uuf__._1363_/X __dut__.__uuf__._1375_/X __dut__._2325_/B
+ __dut__.__uuf__._1363_/X VGND VGND VPWR VPWR __dut__._2324_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1630_ __dut__._1630_/A1 __dut__._1628_/X __dut__._1629_/X VGND VGND VPWR
+ VPWR __dut__._2873_/D sky130_fd_sc_hd__a21o_4
XFILLER_131_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1561_ __dut__._1565_/A __dut__._2855_/Q VGND VGND VPWR VPWR __dut__._1561_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1492_ __dut__._1374_/Y mp[4] __dut__._1491_/X VGND VGND VPWR VPWR __dut__._1492_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_73_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2113_ __dut__._2325_/A __dut__._2113_/B VGND VGND VPWR VPWR __dut__._2113_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._3093_ __dut__._3093_/CLK __dut__._3093_/D __dut__._2525_/Y VGND VGND VPWR
+ VPWR __dut__._3093_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_33_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2044_ __dut__._2044_/A1 prod[4] __dut__._2043_/X VGND VGND VPWR VPWR __dut__._3079_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1749__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3100__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2946_ __dut__._2961_/CLK __dut__._2946_/D __dut__._2672_/Y VGND VGND VPWR
+ VPWR __dut__._2946_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2877_ __dut__._3109_/CLK __dut__._2877_/D __dut__._2741_/Y VGND VGND VPWR
+ VPWR __dut__._2877_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1828_ __dut__._1830_/A1 tie[66] __dut__._1827_/X VGND VGND VPWR VPWR __dut__._2971_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2230__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_122_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1759_ __dut__._2189_/A __dut__._2936_/Q VGND VGND VPWR VPWR __dut__._1759_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_95_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1659__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_297_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1230_ __dut__.__uuf__._1446_/A VGND VGND VPWR VPWR __dut__.__uuf__._1326_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_113_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1161_ __dut__.__uuf__._1161_/A VGND VGND VPWR VPWR __dut__.__uuf__._1161_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_141_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1092_ __dut__.__uuf__._1088_/X __dut__.__uuf__._1085_/X prod[42]
+ prod[43] __dut__.__uuf__._1082_/X VGND VGND VPWR VPWR __dut__._2466_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_95_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1994_ VGND VGND VPWR VPWR __dut__.__uuf__._1994_/HI tie[1] sky130_fd_sc_hd__conb_1
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2800_ rst VGND VGND VPWR VPWR __dut__._2800_/Y sky130_fd_sc_hd__inv_2
X__dut__._2731_ rst VGND VGND VPWR VPWR __dut__._2731_/Y sky130_fd_sc_hd__inv_2
X__dut__._2662_ rst VGND VGND VPWR VPWR __dut__._2662_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1428_ __dut__.__uuf__._1427_/Y __dut__.__uuf__._1423_/X __dut__.__uuf__._1322_/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._1428_/X sky130_fd_sc_hd__o21a_4
XFILLER_49_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1613_ __dut__._2105_/A __dut__._2868_/Q VGND VGND VPWR VPWR __dut__._1613_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1359_ __dut__.__uuf__._1352_/X __dut__.__uuf__._1358_/X __dut__._2331_/B
+ __dut__.__uuf__._1352_/X VGND VGND VPWR VPWR __dut__._2330_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._2593_ rst VGND VGND VPWR VPWR __dut__._2593_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1544_ __dut__._1374_/Y mp[16] __dut__._1543_/X VGND VGND VPWR VPWR __dut__._1544_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1475_ __dut__._2509_/A __dut__._2835_/Q VGND VGND VPWR VPWR __dut__._1475_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_100_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_2_0___dut__.__uuf__.__clk_source__ clkbuf_4_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2251_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1680__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3076_ __dut__._3079_/CLK __dut__._3076_/D __dut__._2542_/Y VGND VGND VPWR
+ VPWR __dut__._3076_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1432__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2027_ __dut__._2207_/A __dut__._3070_/Q VGND VGND VPWR VPWR __dut__._2027_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_285_ _290_/CLK _285_/D VGND VGND VPWR VPWR _285_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1479__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_7_0___dut__.__uuf__.__clk_source___A clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2929_ clkbuf_5_0_0_tck/X __dut__._2929_/D __dut__._2689_/Y VGND VGND VPWR
+ VPWR __dut__._2929_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_114_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2773__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_212_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2276__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1389__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2331_ __dut__.__uuf__._2358_/CLK __dut__._2442_/X __dut__.__uuf__._1125_/X
+ VGND VGND VPWR VPWR prod[30] sky130_fd_sc_hd__dfrtp_4
XFILLER_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2262_ __dut__.__uuf__._2293_/CLK __dut__._2304_/X __dut__.__uuf__._1421_/X
+ VGND VGND VPWR VPWR __dut__._2305_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1213_ __dut__.__uuf__._1234_/A VGND VGND VPWR VPWR __dut__.__uuf__._1213_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_102_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2013__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2193_ __dut__.__uuf__._2216_/CLK __dut__._2166_/X __dut__.__uuf__._1611_/X
+ VGND VGND VPWR VPWR __dut__._2167_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_113_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1144_ __dut__.__uuf__._1173_/A VGND VGND VPWR VPWR __dut__.__uuf__._1144_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1075_ __dut__.__uuf__._1640_/A VGND VGND VPWR VPWR __dut__.__uuf__._1134_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_83_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1662__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2683__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1977_ __dut__.__uuf__._1970_/A __dut__.__uuf__._1975_/B __dut__.__uuf__._1936_/X
+ VGND VGND VPWR VPWR __dut__._2230_/A2 sky130_fd_sc_hd__o21a_4
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3019__CLK clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_tck clkbuf_0_tck/X VGND VGND VPWR VPWR clkbuf_2_3_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2714_ rst VGND VGND VPWR VPWR __dut__._2714_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2645_ rst VGND VGND VPWR VPWR __dut__._2645_/Y sky130_fd_sc_hd__inv_2
X__dut__._2576_ rst VGND VGND VPWR VPWR __dut__._2576_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1527_ __dut__._2509_/A __dut__._2848_/Q VGND VGND VPWR VPWR __dut__._1527_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1458_ __dut__._1458_/A1 __dut__._1456_/X __dut__._1457_/X VGND VGND VPWR
+ VPWR __dut__._2830_/D sky130_fd_sc_hd__a21o_4
XFILLER_132_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1389_ __dut__._2189_/A __dut__._2812_/Q VGND VGND VPWR VPWR __dut__._1389_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2593__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2299__CLK __dut__.__uuf__._2303_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._3059_ __dut__._3059_/CLK __dut__._3059_/D __dut__._2559_/Y VGND VGND VPWR
+ VPWR __dut__._3059_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_268_ _274_/CLK _268_/D VGND VGND VPWR VPWR _268_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_199_ _199_/A VGND VGND VPWR VPWR _199_/X sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1937__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_psn_inst_psn_buff_162_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2768__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1892__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1644__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1900_ __dut__.__uuf__._1867_/X __dut__.__uuf__._1898_/B __dut__.__uuf__._1898_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1901_/C sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1831_ __dut__._2179_/B __dut__._2185_/B VGND VGND VPWR VPWR __dut__.__uuf__._1832_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_33_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1762_ __dut__.__uuf__._1762_/A VGND VGND VPWR VPWR __dut__._2152_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1693_ __dut__.__uuf__._1261_/X __dut__.__uuf__._1691_/B __dut__.__uuf__._1691_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1694_/C sky130_fd_sc_hd__o21a_4
XFILLER_119_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2314_ __dut__.__uuf__._2358_/CLK __dut__._2408_/X __dut__.__uuf__._1175_/X
+ VGND VGND VPWR VPWR prod[13] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2245_ __dut__.__uuf__._2251_/CLK __dut__._2270_/X __dut__.__uuf__._1498_/X
+ VGND VGND VPWR VPWR __dut__._2271_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2176_ __dut__.__uuf__._2225_/CLK __dut__._2132_/X __dut__.__uuf__._1631_/X
+ VGND VGND VPWR VPWR __dut__._2133_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2430_ __dut__._2430_/A1 __dut__._2430_/A2 __dut__._2429_/X VGND VGND VPWR
+ VPWR __dut__._2430_/X sky130_fd_sc_hd__a21o_4
XFILLER_102_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2678__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1127_ __dut__.__uuf__._1118_/X __dut__.__uuf__._1115_/X prod[30]
+ prod[31] __dut__.__uuf__._1126_/X VGND VGND VPWR VPWR __dut__._2442_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_46_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2397__B prod[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2361_ __dut__._2407_/A __dut__._2361_/B VGND VGND VPWR VPWR __dut__._2361_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_83_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1058_ __dut__.__uuf__._1057_/X __dut__.__uuf__._1054_/X prod[53]
+ prod[54] __dut__.__uuf__._1051_/X VGND VGND VPWR VPWR __dut__._2488_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._2292_ __dut__._2292_/A1 __dut__._2292_/A2 __dut__._2291_/X VGND VGND VPWR
+ VPWR __dut__._2292_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2060__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_122_ _291_/Q VGND VGND VPWR VPWR _231_/A sky130_fd_sc_hd__buf_2
XFILLER_137_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1757__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2628_ rst VGND VGND VPWR VPWR __dut__._2628_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2588__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2559_ rst VGND VGND VPWR VPWR __dut__._2559_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1667__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2030_ VGND VGND VPWR VPWR __dut__.__uuf__._2030_/HI tie[37] sky130_fd_sc_hd__conb_1
XFILLER_111_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_17_0_tck clkbuf_4_8_0_tck/X VGND VGND VPWR VPWR __dut__._3079_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1814_ __dut__.__uuf__._1813_/X __dut__.__uuf__._1811_/B __dut__.__uuf__._1811_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1815_/C sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1745_ __dut__.__uuf__._1745_/A VGND VGND VPWR VPWR __dut__.__uuf__._1745_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1930_ __dut__._1930_/A1 tie[117] __dut__._1929_/X VGND VGND VPWR VPWR __dut__._3022_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_119_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1676_ __dut__._1464_/X VGND VGND VPWR VPWR __dut__.__uuf__._1680_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_106_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1861_ __dut__._1881_/A __dut__._2987_/Q VGND VGND VPWR VPWR __dut__._1861_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1792_ __dut__._1830_/A1 tie[48] __dut__._1791_/X VGND VGND VPWR VPWR __dut__._2953_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__275__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2228_ __dut__.__uuf__._2291_/CLK __dut__._2236_/X __dut__.__uuf__._1567_/X
+ VGND VGND VPWR VPWR __dut__._2237_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2159_ VGND VGND VPWR VPWR __dut__.__uuf__._2159_/HI tie[166] sky130_fd_sc_hd__conb_1
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2413_ __dut__._2415_/A prod[15] VGND VGND VPWR VPWR __dut__._2413_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2201__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1608__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2344_ __dut__._2368_/A1 __dut__._2344_/A2 __dut__._2343_/X VGND VGND VPWR
+ VPWR __dut__._2344_/X sky130_fd_sc_hd__a21o_4
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_63_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2275_ __dut__._2281_/A __dut__._2275_/B VGND VGND VPWR VPWR __dut__._2275_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1487__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._2111__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_125_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1530_ __dut__._1516_/X __dut__.__uuf__._1529_/X __dut__._2259_/B
+ __dut__.__uuf__._1513_/X VGND VGND VPWR VPWR __dut__.__uuf__._1530_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__._2781__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1397__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1461_ __dut__.__uuf__._1461_/A VGND VGND VPWR VPWR __dut__.__uuf__._1479_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_143_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1392_ __dut__.__uuf__._1411_/A VGND VGND VPWR VPWR __dut__.__uuf__._1392_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_0_0_tck clkbuf_5_1_0_tck/A VGND VGND VPWR VPWR clkbuf_5_0_0_tck/X sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._2021__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2013_ VGND VGND VPWR VPWR __dut__.__uuf__._2013_/HI tie[20] sky130_fd_sc_hd__conb_1
XFILLER_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2060_ __dut__._2412_/A1 prod[12] __dut__._2059_/X VGND VGND VPWR VPWR __dut__._3087_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_53_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2691__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1728_ __dut__.__uuf__._1704_/X __dut__.__uuf__._1726_/B __dut__.__uuf__._1726_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1729_/C sky130_fd_sc_hd__o21a_4
X__dut__._2962_ __dut__._3079_/CLK __dut__._2962_/D __dut__._2656_/Y VGND VGND VPWR
+ VPWR __dut__._2962_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1913_ __dut__._2005_/A __dut__._3013_/Q VGND VGND VPWR VPWR __dut__._1913_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1659_ __dut__.__uuf__._1706_/A __dut__.__uuf__._1659_/B __dut__.__uuf__._1659_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1660_/A sky130_fd_sc_hd__or3_4
XFILLER_146_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2893_ __dut__._3106_/CLK __dut__._2893_/D __dut__._2725_/Y VGND VGND VPWR
+ VPWR __dut__._2893_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1844_ __dut__._1844_/A1 tie[74] __dut__._1843_/X VGND VGND VPWR VPWR __dut__._2979_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1775_ __dut__._1775_/A __dut__._2944_/Q VGND VGND VPWR VPWR __dut__._1775_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_103_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2327_ __dut__._2407_/A __dut__._2327_/B VGND VGND VPWR VPWR __dut__._2327_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_44_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2258_ __dut__._2262_/A1 __dut__._2258_/A2 __dut__._2257_/X VGND VGND VPWR
+ VPWR __dut__._2258_/X sky130_fd_sc_hd__a21o_4
XFILLER_16_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_121 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1848_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_110 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1820_/A1 sky130_fd_sc_hd__buf_2
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_132 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1884_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_143 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2434_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2189_ __dut__._2189_/A __dut__._2189_/B VGND VGND VPWR VPWR __dut__._2189_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_154 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2448_/A1 sky130_fd_sc_hd__buf_2
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__314__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_176 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1562_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_187 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._1760_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_198 psn_inst_psn_buff_201/A VGND VGND VPWR VPWR __dut__._2200_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_165 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1688_/A1 sky130_fd_sc_hd__buf_2
XFILLER_129_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1945__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_242_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2776__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2495__B prod[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1513_ __dut__.__uuf__._1709_/A VGND VGND VPWR VPWR __dut__.__uuf__._1513_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_128_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1444_ __dut__.__uuf__._1440_/X __dut__.__uuf__._1435_/X __dut__._2297_/B
+ __dut__.__uuf__._1988_/B __dut__.__uuf__._1443_/X VGND VGND VPWR VPWR __dut__._2296_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_132_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1375_ __dut__.__uuf__._1372_/Y __dut__.__uuf__._1373_/X __dut__.__uuf__._1374_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1375_/X sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._3052__CLK __dut__._3059_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1560_ __dut__._1374_/Y mp[19] __dut__._1559_/X VGND VGND VPWR VPWR __dut__._1560_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1491_ __dut__._2509_/A __dut__._2839_/Q VGND VGND VPWR VPWR __dut__._1491_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2484__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2686__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2182__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._3092_ __dut__._3093_/CLK __dut__._3092_/D __dut__._2526_/Y VGND VGND VPWR
+ VPWR __dut__._3092_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2112_ __dut__._2112_/A1 __dut__._2112_/A2 __dut__._2111_/X VGND VGND VPWR
+ VPWR __dut__._2112_/X sky130_fd_sc_hd__a21o_4
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2043_ __dut__._2389_/A __dut__._3078_/Q VGND VGND VPWR VPWR __dut__._2043_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_22_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_26_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2945_ __dut__._2958_/CLK __dut__._2945_/D __dut__._2673_/Y VGND VGND VPWR
+ VPWR __dut__._2945_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_7_0_tck clkbuf_4_7_0_tck/A VGND VGND VPWR VPWR clkbuf_4_7_0_tck/X sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__.__uuf__._1031__B1 prod[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2876_ __dut__._3109_/CLK __dut__._2876_/D __dut__._2742_/Y VGND VGND VPWR
+ VPWR __dut__._2876_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1827_ __dut__._2507_/A __dut__._2970_/Q VGND VGND VPWR VPWR __dut__._1827_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_79_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1758_ __dut__._1760_/A1 tie[31] __dut__._1757_/X VGND VGND VPWR VPWR __dut__._2936_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA_clkbuf_3_2_0___dut__.__uuf__.__clk_source___A clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1689_ __dut__._1689_/A __dut__._2901_/Q VGND VGND VPWR VPWR __dut__._1689_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2596__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3075__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1675__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1160_ __dut__.__uuf__._1147_/X __dut__.__uuf__._1159_/X prod[19]
+ prod[20] __dut__.__uuf__._1156_/X VGND VGND VPWR VPWR __dut__._2420_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2466__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1091_ __dut__.__uuf__._1101_/A VGND VGND VPWR VPWR __dut__.__uuf__._1091_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_67_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1993_ VGND VGND VPWR VPWR __dut__.__uuf__._1993_/HI tie[0] sky130_fd_sc_hd__conb_1
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2730_ rst VGND VGND VPWR VPWR __dut__._2730_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2661_ rst VGND VGND VPWR VPWR __dut__._2661_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1427_ __dut__._2305_/B VGND VGND VPWR VPWR __dut__.__uuf__._1427_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1358_ __dut__.__uuf__._1357_/Y __dut__.__uuf__._1347_/X __dut__.__uuf__._1348_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1358_/X sky130_fd_sc_hd__o21a_4
X__dut__._1612_ __dut__._1374_/Y mp[31] __dut__._1611_/X VGND VGND VPWR VPWR __dut__._1612_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._1564__B2 __dut__.__uuf__._1294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2592_ rst VGND VGND VPWR VPWR __dut__._2592_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1543_ __dut__._2509_/A __dut__._2852_/Q VGND VGND VPWR VPWR __dut__._1543_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1289_ __dut__.__uuf__._1283_/X __dut__.__uuf__._1288_/X __dut__._2357_/B
+ __dut__.__uuf__._1283_/X VGND VGND VPWR VPWR __dut__._2356_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1474_ __dut__._1474_/A1 __dut__._1472_/X __dut__._1473_/X VGND VGND VPWR
+ VPWR __dut__._2834_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1680__A2 prod[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3075_ __dut__._3093_/CLK __dut__._3075_/D __dut__._2543_/Y VGND VGND VPWR
+ VPWR __dut__._3075_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1432__A2 mc[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2026_ __dut__._2026_/A1 tie[165] __dut__._2025_/X VGND VGND VPWR VPWR __dut__._3070_/D
+ sky130_fd_sc_hd__a21o_4
X_284_ _290_/CLK _284_/D VGND VGND VPWR VPWR _284_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._3098__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2928_ clkbuf_5_0_0_tck/X __dut__._2928_/D __dut__._2690_/Y VGND VGND VPWR
+ VPWR __dut__._2928_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1495__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2859_ __dut__._2961_/CLK __dut__._2859_/D __dut__._2759_/Y VGND VGND VPWR
+ VPWR __dut__._2859_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2935__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_205_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_12_0___dut__.__uuf__.__clk_source__ clkbuf_3_6_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2307_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2330_ __dut__.__uuf__._2358_/CLK __dut__._2440_/X __dut__.__uuf__._1128_/X
+ VGND VGND VPWR VPWR prod[29] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2261_ __dut__.__uuf__._2293_/CLK __dut__._2302_/X __dut__.__uuf__._1426_/X
+ VGND VGND VPWR VPWR __dut__._2303_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_114_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1212_ __dut__.__uuf__._1206_/X __dut__.__uuf__._1203_/X prod[1]
+ prod[2] __dut__.__uuf__._1200_/X VGND VGND VPWR VPWR __dut__._2384_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_102_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2192_ __dut__.__uuf__._2216_/CLK __dut__._2164_/X __dut__.__uuf__._1612_/X
+ VGND VGND VPWR VPWR __dut__._2165_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_113_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1143_ __dut__.__uuf__._1146_/A VGND VGND VPWR VPWR __dut__.__uuf__._1143_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_142_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1074_ __dut__.__uuf__._1074_/A VGND VGND VPWR VPWR __dut__.__uuf__._1640_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1976_ __dut__.__uuf__._1976_/A VGND VGND VPWR VPWR __dut__._2232_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_143_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2713_ rst VGND VGND VPWR VPWR __dut__._2713_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2644_ rst VGND VGND VPWR VPWR __dut__._2644_/Y sky130_fd_sc_hd__inv_2
X__dut__._2575_ rst VGND VGND VPWR VPWR __dut__._2575_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_93_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1526_ __dut__._1526_/A1 __dut__._1524_/X __dut__._1525_/X VGND VGND VPWR
+ VPWR __dut__._2847_/D sky130_fd_sc_hd__a21o_4
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1457_ __dut__._2325_/A __dut__._2829_/Q VGND VGND VPWR VPWR __dut__._1457_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1388_ __dut__._1374_/Y mc[12] __dut__._1387_/X VGND VGND VPWR VPWR __dut__._1388_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._3058_ __dut__._3058_/CLK __dut__._3058_/D __dut__._2560_/Y VGND VGND VPWR
+ VPWR __dut__._3058_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._2009_ __dut__._2207_/A __dut__._3061_/Q VGND VGND VPWR VPWR __dut__._2009_/X
+ sky130_fd_sc_hd__and2_4
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_267_ _194_/A _267_/D VGND VGND VPWR VPWR _267_/Q sky130_fd_sc_hd__dfxtp_4
X_198_ _199_/A VGND VGND VPWR VPWR _198_/X sky130_fd_sc_hd__buf_2
XFILLER_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1953__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_155_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2784__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1830_ __dut__._1404_/X VGND VGND VPWR VPWR __dut__.__uuf__._1834_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1761_ __dut__.__uuf__._1761_/A __dut__.__uuf__._1761_/B __dut__.__uuf__._1761_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1762_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1692_ __dut__.__uuf__._1692_/A VGND VGND VPWR VPWR __dut__.__uuf__._1694_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_146_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1580__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2313_ __dut__.__uuf__._2334_/CLK __dut__._2406_/X __dut__.__uuf__._1180_/X
+ VGND VGND VPWR VPWR prod[12] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2244_ __dut__.__uuf__._2251_/CLK __dut__._2268_/X __dut__.__uuf__._1501_/X
+ VGND VGND VPWR VPWR __dut__._2269_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2175_ __dut__.__uuf__._2225_/CLK __dut__._2130_/X __dut__.__uuf__._1632_/X
+ VGND VGND VPWR VPWR __dut__._2131_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1126_ __dut__.__uuf__._1126_/A VGND VGND VPWR VPWR __dut__.__uuf__._1126_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2360_ __dut__._2368_/A1 __dut__._2360_/A2 __dut__._2359_/X VGND VGND VPWR
+ VPWR __dut__._2360_/X sky130_fd_sc_hd__a21o_4
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1057_ __dut__.__uuf__._1088_/A VGND VGND VPWR VPWR __dut__.__uuf__._1057_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2291_ __dut__._2303_/A __dut__._2291_/B VGND VGND VPWR VPWR __dut__._2291_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_83_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2694__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2060__A2 prod[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1959_ __dut__._2227_/B __dut__._2233_/B VGND VGND VPWR VPWR __dut__.__uuf__._1960_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_121_ _310_/Q VGND VGND VPWR VPWR _121_/Y sky130_fd_sc_hd__inv_2
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2627_ rst VGND VGND VPWR VPWR __dut__._2627_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2558_ rst VGND VGND VPWR VPWR __dut__._2558_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2266__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2489_ __dut__._2491_/A prod[53] VGND VGND VPWR VPWR __dut__._2489_/X sky130_fd_sc_hd__and2_4
X__dut__._1509_ __dut__._1509_/A __dut__._2832_/Q VGND VGND VPWR VPWR __dut__._1509_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_19_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2109__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_272_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2779__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._3009__CLK _274_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0_0_tck clkbuf_0_tck/X VGND VGND VPWR VPWR clkbuf_2_1_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._2019__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1813_ __dut__.__uuf__._1921_/A VGND VGND VPWR VPWR __dut__.__uuf__._1813_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1744_ __dut__._2147_/B __dut__._2153_/B VGND VGND VPWR VPWR __dut__.__uuf__._1745_/A
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1675_ __dut__.__uuf__._1668_/A __dut__.__uuf__._1673_/B __dut__.__uuf__._1661_/X
+ VGND VGND VPWR VPWR __dut__._2118_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_146_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1860_ __dut__._1864_/A1 tie[82] __dut__._1859_/X VGND VGND VPWR VPWR __dut__._2987_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1791_ __dut__._1797_/A __dut__._2952_/Q VGND VGND VPWR VPWR __dut__._1791_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2289__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2689__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2227_ __dut__.__uuf__._2291_/CLK __dut__._2234_/X __dut__.__uuf__._1568_/X
+ VGND VGND VPWR VPWR __dut__._2235_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_130_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2158_ VGND VGND VPWR VPWR __dut__.__uuf__._2158_/HI tie[165] sky130_fd_sc_hd__conb_1
X__dut__._2412_ __dut__._2412_/A1 __dut__._2412_/A2 __dut__._2411_/X VGND VGND VPWR
+ VPWR __dut__._2412_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2089_ VGND VGND VPWR VPWR __dut__.__uuf__._2089_/HI tie[96] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1109_ __dut__.__uuf__._1103_/X __dut__.__uuf__._1099_/X prod[36]
+ prod[37] __dut__.__uuf__._1096_/X VGND VGND VPWR VPWR __dut__._2454_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._2343_ __dut__._2407_/A __dut__._2343_/B VGND VGND VPWR VPWR __dut__._2343_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1608__A2 mp[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2274_ __dut__._2278_/A1 __dut__._2274_/A2 __dut__._2273_/X VGND VGND VPWR
+ VPWR __dut__._2274_/X sky130_fd_sc_hd__a21o_4
XFILLER_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1544__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1989_ __dut__._2005_/A __dut__._3051_/Q VGND VGND VPWR VPWR __dut__._1989_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2599__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_psn_inst_psn_buff_118_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1460_ __dut__.__uuf__._1440_/X __dut__.__uuf__._1458_/X __dut__._2289_/B
+ __dut__.__uuf__._1447_/X __dut__.__uuf__._1459_/X VGND VGND VPWR VPWR __dut__._2288_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_155_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1391_ __dut__.__uuf__._1461_/A VGND VGND VPWR VPWR __dut__.__uuf__._1411_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_131_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2012_ VGND VGND VPWR VPWR __dut__.__uuf__._2012_/HI tie[19] sky130_fd_sc_hd__conb_1
XFILLER_150_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1727_ __dut__.__uuf__._1727_/A VGND VGND VPWR VPWR __dut__.__uuf__._1729_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._2961_ __dut__._2961_/CLK __dut__._2961_/D __dut__._2657_/Y VGND VGND VPWR
+ VPWR __dut__._2961_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1912_ __dut__._2004_/A1 tie[108] __dut__._1911_/X VGND VGND VPWR VPWR __dut__._3013_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2892_ __dut__._3102_/CLK __dut__._2892_/D __dut__._2726_/Y VGND VGND VPWR
+ VPWR __dut__._2892_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1658_ __dut__.__uuf__._1261_/X __dut__.__uuf__._1656_/B __dut__.__uuf__._1656_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1659_/C sky130_fd_sc_hd__o21a_4
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1843_ __dut__._1843_/A __dut__._2978_/Q VGND VGND VPWR VPWR __dut__._1843_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1589_ __dut__.__uuf__._1590_/A VGND VGND VPWR VPWR __dut__.__uuf__._1589_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1774_ __dut__._1780_/A1 tie[39] __dut__._1773_/X VGND VGND VPWR VPWR __dut__._2944_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2326_ __dut__._2332_/A1 __dut__._2326_/A2 __dut__._2325_/X VGND VGND VPWR
+ VPWR __dut__._2326_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2257_ __dut__._2257_/A __dut__._2257_/B VGND VGND VPWR VPWR __dut__._2257_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_111 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1830_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_100 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1780_/A1 sky130_fd_sc_hd__buf_4
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_122 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1864_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_133 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1886_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_144 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2436_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2188_ __dut__._2192_/A1 __dut__._2188_/A2 __dut__._2187_/X VGND VGND VPWR
+ VPWR __dut__._2188_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_155 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2098_/A1 sky130_fd_sc_hd__buf_2
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_177 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2256_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_188 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._1942_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_166 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2504_/A1 sky130_fd_sc_hd__buf_2
XFILLER_129_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_16_0_tck clkbuf_4_8_0_tck/X VGND VGND VPWR VPWR __dut__._2985_/CLK sky130_fd_sc_hd__clkbuf_1
Xpsn_inst_psn_buff_199 psn_inst_psn_buff_201/A VGND VGND VPWR VPWR __dut__._2208_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_144_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1961__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_235_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2792__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1512_ __dut__.__uuf__._1533_/A VGND VGND VPWR VPWR __dut__.__uuf__._1512_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1443_ __dut__._1604_/X __dut__.__uuf__._1442_/X __dut__._2299_/B
+ __dut__.__uuf__._1423_/X VGND VGND VPWR VPWR __dut__.__uuf__._1443_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__._1508__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1374_ __dut__.__uuf__._1399_/A VGND VGND VPWR VPWR __dut__.__uuf__._1374_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2991__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1490_ __dut__._1490_/A1 __dut__._1488_/X __dut__._1489_/X VGND VGND VPWR
+ VPWR __dut__._2838_/D sky130_fd_sc_hd__a21o_4
XFILLER_100_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3091_ __dut__._3093_/CLK __dut__._3091_/D __dut__._2527_/Y VGND VGND VPWR
+ VPWR __dut__._3091_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2111_ __dut__._2325_/A __dut__._2111_/B VGND VGND VPWR VPWR __dut__._2111_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2042_ __dut__._2044_/A1 prod[3] __dut__._2041_/X VGND VGND VPWR VPWR __dut__._3078_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_110_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2207__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_19_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2944_ __dut__._2958_/CLK __dut__._2944_/D __dut__._2674_/Y VGND VGND VPWR
+ VPWR __dut__._2944_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1031__B2 __dut__.__uuf__._1025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2875_ __dut__._3109_/CLK __dut__._2875_/D __dut__._2743_/Y VGND VGND VPWR
+ VPWR __dut__._2875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1826_ __dut__._1830_/A1 tie[65] __dut__._1825_/X VGND VGND VPWR VPWR __dut__._2970_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2172__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1757_ __dut__._2189_/A __dut__._2935_/Q VGND VGND VPWR VPWR __dut__._1757_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1688_ __dut__._1688_/A1 prod[61] __dut__._1687_/X VGND VGND VPWR VPWR __dut__._2901_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_95_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2309_ __dut__._2325_/A __dut__._2309_/B VGND VGND VPWR VPWR __dut__._2309_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1986__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__288__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2117__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1910__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1090_ __dut__.__uuf__._1134_/A VGND VGND VPWR VPWR __dut__.__uuf__._1101_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2787__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1691__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1992_ __dut__.__uuf__._1992_/A VGND VGND VPWR VPWR __dut__.__uuf__._1992_/X
+ sky130_fd_sc_hd__buf_2
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2027__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2154__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2660_ rst VGND VGND VPWR VPWR __dut__._2660_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1426_ __dut__.__uuf__._1434_/A VGND VGND VPWR VPWR __dut__.__uuf__._1426_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1357_ __dut__._2333_/B VGND VGND VPWR VPWR __dut__.__uuf__._1357_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1611_ __dut__._2509_/A __dut__._2869_/Q VGND VGND VPWR VPWR __dut__._1611_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2591_ rst VGND VGND VPWR VPWR __dut__._2591_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2697__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1542_ __dut__._1562_/A1 __dut__._1540_/X __dut__._1541_/X VGND VGND VPWR
+ VPWR __dut__._2851_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1288_ __dut__.__uuf__._1287_/Y __dut__.__uuf__._1985_/A __dut__.__uuf__._1268_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1288_/X sky130_fd_sc_hd__o21a_4
XFILLER_46_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1473_ __dut__._2281_/A __dut__._2833_/Q VGND VGND VPWR VPWR __dut__._1473_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_105_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2887__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3074_ _194_/A __dut__._3074_/D __dut__._2544_/Y VGND VGND VPWR VPWR _210_/A2
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1968__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2025_ __dut__._2207_/A __dut__._3069_/Q VGND VGND VPWR VPWR __dut__._2025_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_283_ _290_/CLK _283_/D VGND VGND VPWR VPWR _283_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2927_ clkbuf_5_9_0_tck/X __dut__._2927_/D __dut__._2691_/Y VGND VGND VPWR
+ VPWR __dut__._2927_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2858_ __dut__._2961_/CLK __dut__._2858_/D __dut__._2760_/Y VGND VGND VPWR
+ VPWR __dut__._2858_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1809_ __dut__._1817_/A __dut__._2961_/Q VGND VGND VPWR VPWR __dut__._1809_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2789_ rst VGND VGND VPWR VPWR __dut__._2789_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3042__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_100_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_9_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._2384__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2172__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2260_ __dut__.__uuf__._2293_/CLK __dut__._2300_/X __dut__.__uuf__._1430_/X
+ VGND VGND VPWR VPWR __dut__._2301_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_141_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1211_ __dut__.__uuf__._1234_/A VGND VGND VPWR VPWR __dut__.__uuf__._1211_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2191_ __dut__.__uuf__._2216_/CLK __dut__._2162_/X __dut__.__uuf__._1613_/X
+ VGND VGND VPWR VPWR __dut__._2163_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1142_ __dut__.__uuf__._1132_/X __dut__.__uuf__._1129_/X prod[25]
+ prod[26] __dut__.__uuf__._1141_/X VGND VGND VPWR VPWR __dut__._2432_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1073_ __dut__.__uuf__._1072_/X __dut__.__uuf__._1069_/X prod[48]
+ prod[49] __dut__.__uuf__._1066_/X VGND VGND VPWR VPWR __dut__._2478_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_83_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_6_0_tck clkbuf_4_7_0_tck/A VGND VGND VPWR VPWR clkbuf_4_6_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1975_ __dut__.__uuf__._1975_/A __dut__.__uuf__._1975_/B __dut__.__uuf__._1975_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1976_/A sky130_fd_sc_hd__or3_4
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2712_ rst VGND VGND VPWR VPWR __dut__._2712_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1409_ __dut__.__uuf__._1408_/Y __dut__.__uuf__._1398_/X __dut__.__uuf__._1399_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1409_/X sky130_fd_sc_hd__o21a_4
X__dut__._2643_ rst VGND VGND VPWR VPWR __dut__._2643_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2574_ rst VGND VGND VPWR VPWR __dut__._2574_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_86_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1525_ __dut__._1557_/A __dut__._2846_/Q VGND VGND VPWR VPWR __dut__._1525_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_86_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1456_ __dut__._1374_/Y mc[28] __dut__._1455_/X VGND VGND VPWR VPWR __dut__._1456_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._3065__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1387_ __dut__._2509_/A __dut__._2813_/Q VGND VGND VPWR VPWR __dut__._1387_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._3057_ _271_/CLK __dut__._3057_/D __dut__._2561_/Y VGND VGND VPWR VPWR __dut__._3057_/Q
+ sky130_fd_sc_hd__dfrtp_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2008_ __dut__._2008_/A1 tie[156] __dut__._2007_/X VGND VGND VPWR VPWR __dut__._3061_/D
+ sky130_fd_sc_hd__a21o_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_266_ _274_/CLK _266_/D VGND VGND VPWR VPWR _266_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__.__uuf__._2195__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2366__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_197_ _199_/A VGND VGND VPWR VPWR _197_/X sky130_fd_sc_hd__buf_2
XFILLER_10_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2902__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_148_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1760_ __dut__.__uuf__._1759_/X __dut__.__uuf__._1757_/B __dut__.__uuf__._1757_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1761_/C sky130_fd_sc_hd__o21a_4
XFILLER_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1691_ __dut__.__uuf__._1736_/A __dut__.__uuf__._1691_/B __dut__.__uuf__._1691_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1692_/A sky130_fd_sc_hd__or3_4
XFILLER_20_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2312_ __dut__.__uuf__._2334_/CLK __dut__._2404_/X __dut__.__uuf__._1182_/X
+ VGND VGND VPWR VPWR prod[11] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2305__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1580__A2 mp[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2243_ __dut__.__uuf__._2251_/CLK __dut__._2266_/X __dut__.__uuf__._1506_/X
+ VGND VGND VPWR VPWR __dut__._2267_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_153_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2174_ __dut__.__uuf__._2225_/CLK __dut__._2128_/X __dut__.__uuf__._1633_/X
+ VGND VGND VPWR VPWR __dut__._2129_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1125_ __dut__.__uuf__._1131_/A VGND VGND VPWR VPWR __dut__.__uuf__._1125_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_68_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3088__CLK __dut__._3106_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1056_ __dut__.__uuf__._1056_/A VGND VGND VPWR VPWR __dut__.__uuf__._1056_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2290_ __dut__._2290_/A1 __dut__._2290_/A2 __dut__._2289_/X VGND VGND VPWR
+ VPWR __dut__._2290_/X sky130_fd_sc_hd__a21o_4
XFILLER_83_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__291__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2925__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1958_ __dut__._1456_/X VGND VGND VPWR VPWR __dut__.__uuf__._1962_/B
+ sky130_fd_sc_hd__inv_2
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1207__A1 __dut__.__uuf__._1206_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1889_ __dut__.__uuf__._1889_/A VGND VGND VPWR VPWR __dut__.__uuf__._1891_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2348__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2215__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2626_ rst VGND VGND VPWR VPWR __dut__._2626_/Y sky130_fd_sc_hd__inv_2
X__dut__._2557_ rst VGND VGND VPWR VPWR __dut__._2557_/Y sky130_fd_sc_hd__inv_2
XANTENNA__308__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2488_ __dut__._2488_/A1 __dut__._2488_/A2 __dut__._2487_/X VGND VGND VPWR
+ VPWR __dut__._2488_/X sky130_fd_sc_hd__a21o_4
X__dut__._1508_ __dut__._1374_/Y mc[3] __dut__._1507_/X VGND VGND VPWR VPWR __dut__._1508_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_62_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1439_ __dut__._2509_/A __dut__._2826_/Q VGND VGND VPWR VPWR __dut__._1439_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_61_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3109_ __dut__._3109_/CLK __dut__._3109_/D __dut__._2809_/Y VGND VGND VPWR
+ VPWR __dut__._3109_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2109__B __dut__._2109_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_249_ _200_/X _313_/Q VGND VGND VPWR VPWR _249_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_143_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2125__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_265_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__.__uuf__._2210__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_111_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2795__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1437__A1 __dut__.__uuf__._1206_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1812_ __dut__.__uuf__._1812_/A VGND VGND VPWR VPWR __dut__.__uuf__._1815_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_61_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1743_ __dut__._1628_/X VGND VGND VPWR VPWR __dut__.__uuf__._1747_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_33_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1674_ __dut__.__uuf__._1674_/A VGND VGND VPWR VPWR __dut__._2120_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1790_ __dut__._1790_/A1 tie[47] __dut__._1789_/X VGND VGND VPWR VPWR __dut__._2952_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2502__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2226_ __dut__.__uuf__._2291_/CLK __dut__._2232_/X __dut__.__uuf__._1569_/X
+ VGND VGND VPWR VPWR __dut__._2233_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_88_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2411_ __dut__._2415_/A prod[14] VGND VGND VPWR VPWR __dut__._2411_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._2157_ VGND VGND VPWR VPWR __dut__.__uuf__._2157_/HI tie[164] sky130_fd_sc_hd__conb_1
XFILLER_76_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2342_ __dut__._2368_/A1 __dut__._2342_/A2 __dut__._2341_/X VGND VGND VPWR
+ VPWR __dut__._2342_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2088_ VGND VGND VPWR VPWR __dut__.__uuf__._2088_/HI tie[95] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1108_ __dut__.__uuf__._1117_/A VGND VGND VPWR VPWR __dut__.__uuf__._1108_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_44_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1039_ __dut__.__uuf__._1464_/A VGND VGND VPWR VPWR __dut__.__uuf__._1099_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._2273_ __dut__._2281_/A __dut__._2273_/B VGND VGND VPWR VPWR __dut__._2273_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_113_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._3103__CLK __dut__._3106_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1544__A2 mp[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2233__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1988_ __dut__._1990_/A1 tie[146] __dut__._1987_/X VGND VGND VPWR VPWR __dut__._3051_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_113_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2609_ rst VGND VGND VPWR VPWR __dut__._2609_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1116__B1 prod[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1480__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1959__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1198__A3 prod[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1390_ __dut__.__uuf__._1378_/X __dut__.__uuf__._1388_/X __dut__._2319_/B
+ __dut__.__uuf__._1389_/X VGND VGND VPWR VPWR __dut__._2318_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2011_ VGND VGND VPWR VPWR __dut__.__uuf__._2011_/HI tie[18] sky130_fd_sc_hd__conb_1
XFILLER_85_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1658__A1 __dut__.__uuf__._1261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1122__A3 prod[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1726_ __dut__.__uuf__._1736_/A __dut__.__uuf__._1726_/B __dut__.__uuf__._1726_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1727_/A sky130_fd_sc_hd__or3_4
X__dut__._2960_ __dut__._2961_/CLK __dut__._2960_/D __dut__._2658_/Y VGND VGND VPWR
+ VPWR __dut__._2960_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1911_ __dut__._2005_/A __dut__._3012_/Q VGND VGND VPWR VPWR __dut__._1911_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2891_ __dut__._3102_/CLK __dut__._2891_/D __dut__._2727_/Y VGND VGND VPWR
+ VPWR __dut__._2891_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1657_ __dut__.__uuf__._1657_/A VGND VGND VPWR VPWR __dut__.__uuf__._1659_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._1842_ __dut__._1842_/A1 tie[73] __dut__._1841_/X VGND VGND VPWR VPWR __dut__._2978_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1588_ __dut__.__uuf__._1590_/A VGND VGND VPWR VPWR __dut__.__uuf__._1588_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1773_ __dut__._1775_/A __dut__._2943_/Q VGND VGND VPWR VPWR __dut__._1773_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2209_ __dut__.__uuf__._2230_/CLK __dut__._2198_/X __dut__.__uuf__._1590_/X
+ VGND VGND VPWR VPWR __dut__._2199_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_130_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2325_ __dut__._2325_/A __dut__._2325_/B VGND VGND VPWR VPWR __dut__._2325_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2256_ __dut__._2256_/A1 __dut__._2256_/A2 __dut__._2255_/X VGND VGND VPWR
+ VPWR __dut__._2256_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_112 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1832_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_101 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1782_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2187_ __dut__._2197_/A __dut__._2187_/B VGND VGND VPWR VPWR __dut__._2187_/X
+ sky130_fd_sc_hd__and2_4
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_123 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1868_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_134 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2078_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_145 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2438_/A1 sky130_fd_sc_hd__buf_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_189 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._2184_/A1
+ sky130_fd_sc_hd__buf_4
Xpsn_inst_psn_buff_178 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR psn_inst_psn_buff_190/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_156 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2100_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_167 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1686_/A1 sky130_fd_sc_hd__buf_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2403__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1961__B __dut__._3037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_130_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_228_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1511_ __dut__.__uuf__._1522_/A VGND VGND VPWR VPWR __dut__.__uuf__._1511_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1114__A __dut__.__uuf__._1464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1442_ __dut__.__uuf__._1563_/A VGND VGND VPWR VPWR __dut__.__uuf__._1442_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1508__A2 mc[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1373_ __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR __dut__.__uuf__._1373_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2313__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1692__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3090_ __dut__._3093_/CLK __dut__._3090_/D __dut__._2528_/Y VGND VGND VPWR
+ VPWR __dut__._3090_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1444__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2110_ __dut__._2110_/A1 __dut__._2110_/A2 __dut__._2109_/X VGND VGND VPWR
+ VPWR __dut__._2110_/X sky130_fd_sc_hd__a21o_4
XFILLER_81_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2041_ __dut__._2041_/A __dut__._3077_/Q VGND VGND VPWR VPWR __dut__._2041_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_14_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1599__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2943_ __dut__._2958_/CLK __dut__._2943_/D __dut__._2675_/Y VGND VGND VPWR
+ VPWR __dut__._2943_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1024__A __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1709_ __dut__.__uuf__._1709_/A VGND VGND VPWR VPWR __dut__.__uuf__._1926_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_126_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2874_ clkbuf_5_2_0_tck/X __dut__._2874_/D __dut__._2744_/Y VGND VGND VPWR
+ VPWR __dut__._2874_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1031__A2 __dut__.__uuf__._1023_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1825_ __dut__._1825_/A __dut__._2969_/Q VGND VGND VPWR VPWR __dut__._1825_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2223__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1756_ __dut__._1760_/A1 tie[30] __dut__._1755_/X VGND VGND VPWR VPWR __dut__._2935_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_135_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1687_ __dut__._1689_/A __dut__._2900_/Q VGND VGND VPWR VPWR __dut__._1687_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_2_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2308_ __dut__._2308_/A1 __dut__._2308_/A2 __dut__._2307_/X VGND VGND VPWR
+ VPWR __dut__._2308_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2239_ __dut__._2245_/A __dut__._2239_/B VGND VGND VPWR VPWR __dut__._2239_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_178_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1264__A1_N __dut__.__uuf__._1261_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_140_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1674__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1991_ done __dut__.__uuf__._1990_/Y __dut__._1616_/X VGND VGND VPWR
+ VPWR __dut__._2108_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_63_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1425_ __dut__.__uuf__._1414_/X __dut__.__uuf__._1424_/X __dut__._2305_/B
+ __dut__.__uuf__._1414_/X VGND VGND VPWR VPWR __dut__._2304_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1356_ __dut__.__uuf__._1360_/A VGND VGND VPWR VPWR __dut__.__uuf__._1356_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1610_ __dut__._1610_/A1 __dut__._1608_/X __dut__._1609_/X VGND VGND VPWR
+ VPWR __dut__._2868_/D sky130_fd_sc_hd__a21o_4
XFILLER_132_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2590_ rst VGND VGND VPWR VPWR __dut__._2590_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1541_ __dut__._1557_/A __dut__._2850_/Q VGND VGND VPWR VPWR __dut__._1541_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1287_ __dut__._2359_/B VGND VGND VPWR VPWR __dut__.__uuf__._1287_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_86_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1472_ __dut__._1374_/Y mc[31] __dut__._1471_/X VGND VGND VPWR VPWR __dut__._1472_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_105_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_15_0_tck clkbuf_4_7_0_tck/X VGND VGND VPWR VPWR __dut__._2961_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_42_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3073_ clkbuf_5_5_0_tck/X __dut__._3073_/D __dut__._2545_/Y VGND VGND VPWR
+ VPWR __dut__._3073_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_121_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2090__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2024_ __dut__._2024_/A1 tie[164] __dut__._2023_/X VGND VGND VPWR VPWR __dut__._3069_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_139_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_282_ _290_/CLK _282_/D VGND VGND VPWR VPWR _282_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_psn_inst_psn_buff_31_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2926_ clkbuf_5_9_0_tck/X __dut__._2926_/D __dut__._2692_/Y VGND VGND VPWR
+ VPWR __dut__._2926_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2857_ __dut__._2860_/CLK __dut__._2857_/D __dut__._2761_/Y VGND VGND VPWR
+ VPWR __dut__._2857_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1808_ __dut__._1816_/A1 tie[56] __dut__._1807_/X VGND VGND VPWR VPWR __dut__._2961_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2788_ rst VGND VGND VPWR VPWR __dut__._2788_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1739_ __dut__._2189_/A __dut__._2926_/Q VGND VGND VPWR VPWR __dut__._1739_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1656__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1408__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_295_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1210_ __dut__.__uuf__._1206_/X __dut__.__uuf__._1203_/X prod[2]
+ prod[3] __dut__.__uuf__._1200_/X VGND VGND VPWR VPWR __dut__._2386_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._2190_ __dut__.__uuf__._2216_/CLK __dut__._2160_/X __dut__.__uuf__._1614_/X
+ VGND VGND VPWR VPWR __dut__._2161_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_141_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2798__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1141_ __dut__.__uuf__._1200_/A VGND VGND VPWR VPWR __dut__.__uuf__._1141_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1072_ __dut__.__uuf__._1088_/A VGND VGND VPWR VPWR __dut__.__uuf__._1072_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1974_ __dut__.__uuf__._1680_/A __dut__.__uuf__._1972_/B __dut__.__uuf__._1972_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1975_/C sky130_fd_sc_hd__o21a_4
XFILLER_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2711_ rst VGND VGND VPWR VPWR __dut__._2711_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1408_ __dut__._2313_/B VGND VGND VPWR VPWR __dut__.__uuf__._1408_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_116_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2642_ rst VGND VGND VPWR VPWR __dut__._2642_/Y sky130_fd_sc_hd__inv_2
X__dut__._2573_ rst VGND VGND VPWR VPWR __dut__._2573_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1339_ __dut__.__uuf__._1327_/X __dut__.__uuf__._1337_/X __dut__._2339_/B
+ __dut__.__uuf__._1338_/X VGND VGND VPWR VPWR __dut__._2338_/A2 sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._2854__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1524_ __dut__._1374_/Y mp[11] __dut__._1523_/X VGND VGND VPWR VPWR __dut__._1524_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_79_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__306__SET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1455_ __dut__._2509_/A __dut__._2830_/Q VGND VGND VPWR VPWR __dut__._1455_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1972__A __dut__.__uuf__._1982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1386_ __dut__._1714_/A1 __dut__._1384_/X __dut__._1385_/X VGND VGND VPWR
+ VPWR __dut__._2812_/D sky130_fd_sc_hd__a21o_4
XFILLER_92_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3056_ __dut__._3059_/CLK __dut__._3056_/D __dut__._2562_/Y VGND VGND VPWR
+ VPWR __dut__._3056_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2007_ __dut__._2207_/A __dut__._3060_/Q VGND VGND VPWR VPWR __dut__._2007_/X
+ sky130_fd_sc_hd__and2_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_265_ _194_/A _265_/D VGND VGND VPWR VPWR _265_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_196_ _199_/A VGND VGND VPWR VPWR _196_/X sky130_fd_sc_hd__buf_2
XFILLER_108_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2909_ clkbuf_5_2_0_tck/X __dut__._2909_/D __dut__._2709_/Y VGND VGND VPWR
+ VPWR __dut__._2909_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_142_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1882__A __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2054__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_210_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1690_ __dut__._2127_/B __dut__._2133_/B __dut__.__uuf__._1689_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1691_/C sky130_fd_sc_hd__o21ai_4
XFILLER_20_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1697__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2311_ __dut__.__uuf__._2334_/CLK __dut__._2402_/X __dut__.__uuf__._1184_/X
+ VGND VGND VPWR VPWR prod[10] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2242_ __dut__.__uuf__._2251_/CLK __dut__._2264_/X __dut__.__uuf__._1511_/X
+ VGND VGND VPWR VPWR __dut__._2265_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2877__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2321__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2173_ __dut__.__uuf__._2225_/CLK __dut__._2126_/X __dut__.__uuf__._1635_/X
+ VGND VGND VPWR VPWR __dut__._2127_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1124_ __dut__.__uuf__._1118_/X __dut__.__uuf__._1115_/X prod[31]
+ prod[32] __dut__.__uuf__._1111_/X VGND VGND VPWR VPWR __dut__._2444_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1055_ __dut__.__uuf__._1043_/X __dut__.__uuf__._1054_/X prod[54]
+ prod[55] __dut__.__uuf__._1051_/X VGND VGND VPWR VPWR __dut__._2490_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1016__B __dut__._2109_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1957_ __dut__.__uuf__._1950_/A __dut__.__uuf__._1955_/B __dut__.__uuf__._1936_/X
+ VGND VGND VPWR VPWR __dut__._2222_/A2 sky130_fd_sc_hd__o21a_4
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1888_ __dut__.__uuf__._1898_/A __dut__.__uuf__._1888_/B __dut__.__uuf__._1888_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1889_/A sky130_fd_sc_hd__or3_4
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2625_ rst VGND VGND VPWR VPWR __dut__._2625_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2231__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3032__CLK clkbuf_5_1_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2556_ rst VGND VGND VPWR VPWR __dut__._2556_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2487_ __dut__._2491_/A prod[52] VGND VGND VPWR VPWR __dut__._2487_/X sky130_fd_sc_hd__and2_4
X__dut__._1507_ __dut__._2509_/A __dut__._2843_/Q VGND VGND VPWR VPWR __dut__._1507_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_100_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1438_ __dut__._1438_/A1 __dut__._1436_/X __dut__._1437_/X VGND VGND VPWR
+ VPWR __dut__._2825_/D sky130_fd_sc_hd__a21o_4
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3108_ __dut__._3109_/CLK __dut__._3108_/D __dut__._1372_/Y VGND VGND VPWR
+ VPWR __dut__._3108_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._3039_ _306_/CLK __dut__._3039_/D __dut__._2579_/Y VGND VGND VPWR VPWR __dut__._3039_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_156_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_248_ _201_/X _312_/Q VGND VGND VPWR VPWR _248_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_179_ _273_/Q _182_/B VGND VGND VPWR VPWR _272_/D sky130_fd_sc_hd__and2_4
XFILLER_143_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_tck clkbuf_4_5_0_tck/A VGND VGND VPWR VPWR clkbuf_4_5_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_160_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_258_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1811_ __dut__.__uuf__._1844_/A __dut__.__uuf__._1811_/B __dut__.__uuf__._1811_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1812_/A sky130_fd_sc_hd__or3_4
XFILLER_61_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1742_ __dut__.__uuf__._1904_/A VGND VGND VPWR VPWR __dut__.__uuf__._1790_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1673_ __dut__.__uuf__._1706_/A __dut__.__uuf__._1673_/B __dut__.__uuf__._1673_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1674_/A sky130_fd_sc_hd__or3_4
XANTENNA___dut__._2035__B prod[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3055__CLK __dut__._3059_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2051__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2225_ __dut__.__uuf__._2225_/CLK __dut__._2230_/X __dut__.__uuf__._1570_/X
+ VGND VGND VPWR VPWR __dut__._2231_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_130_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2156_ VGND VGND VPWR VPWR __dut__.__uuf__._2156_/HI tie[163] sky130_fd_sc_hd__conb_1
XFILLER_102_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2410_ __dut__._2412_/A1 __dut__._2410_/A2 __dut__._2409_/X VGND VGND VPWR
+ VPWR __dut__._2410_/X sky130_fd_sc_hd__a21o_4
XFILLER_76_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1107_ __dut__.__uuf__._1103_/X __dut__.__uuf__._1099_/X prod[37]
+ prod[38] __dut__.__uuf__._1096_/X VGND VGND VPWR VPWR __dut__._2456_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_113_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2341_ __dut__._2407_/A __dut__._2341_/B VGND VGND VPWR VPWR __dut__._2341_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2185__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2087_ VGND VGND VPWR VPWR __dut__.__uuf__._2087_/HI tie[94] sky130_fd_sc_hd__conb_1
XFILLER_71_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2272_ __dut__._2278_/A1 __dut__._2272_/A2 __dut__._2271_/X VGND VGND VPWR
+ VPWR __dut__._2272_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1038_ __dut__.__uuf__._1042_/A VGND VGND VPWR VPWR __dut__.__uuf__._1038_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_113_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1027__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1987_ __dut__._2005_/A __dut__._3050_/Q VGND VGND VPWR VPWR __dut__._1987_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_125_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2608_ rst VGND VGND VPWR VPWR __dut__._2608_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2539_ rst VGND VGND VPWR VPWR __dut__._2539_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_7_0_tck_A clkbuf_3_7_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1480__A2 mp[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3078__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1052__B1 prod[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1975__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2010_ VGND VGND VPWR VPWR __dut__.__uuf__._2010_/HI tie[17] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2496__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2915__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1725_ __dut__._2139_/B __dut__._2145_/B __dut__.__uuf__._1724_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1726_/C sky130_fd_sc_hd__o21ai_4
XFILLER_119_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1910_ __dut__._2004_/A1 tie[107] __dut__._1909_/X VGND VGND VPWR VPWR __dut__._3012_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1656_ __dut__.__uuf__._1680_/A __dut__.__uuf__._1656_/B __dut__.__uuf__._1656_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1657_/A sky130_fd_sc_hd__or3_4
X__dut__._2890_ __dut__._3102_/CLK __dut__._2890_/D __dut__._2728_/Y VGND VGND VPWR
+ VPWR __dut__._2890_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1841_ __dut__._2507_/A __dut__._2977_/Q VGND VGND VPWR VPWR __dut__._1841_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1587_ __dut__.__uuf__._1590_/A VGND VGND VPWR VPWR __dut__.__uuf__._1587_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_108_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1772_ __dut__._1780_/A1 tie[38] __dut__._1771_/X VGND VGND VPWR VPWR __dut__._2943_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2208_ __dut__.__uuf__._2230_/CLK __dut__._2196_/X __dut__.__uuf__._1592_/X
+ VGND VGND VPWR VPWR __dut__._2197_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2139_ VGND VGND VPWR VPWR __dut__.__uuf__._2139_/HI tie[146] sky130_fd_sc_hd__conb_1
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2324_ __dut__._2332_/A1 __dut__._2324_/A2 __dut__._2323_/X VGND VGND VPWR
+ VPWR __dut__._2324_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_61_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2255_ __dut__._2255_/A __dut__._2255_/B VGND VGND VPWR VPWR __dut__._2255_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpsn_inst_psn_buff_102 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1784_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2186_ __dut__._2192_/A1 __dut__._2186_/A2 __dut__._2185_/X VGND VGND VPWR
+ VPWR __dut__._2186_/X sky130_fd_sc_hd__a21o_4
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_124 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1866_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_113 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1834_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_135 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2076_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_146 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2092_/A1 sky130_fd_sc_hd__buf_2
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__.__uuf__._2200__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_179 psn_inst_psn_buff_190/A VGND VGND VPWR VPWR __dut__._1622_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_157 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2102_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_168 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2502_/A1 sky130_fd_sc_hd__buf_4
XFILLER_40_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2403__B prod[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2478__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_123_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2402__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1510_ __dut__.__uuf__._1507_/X __dut__.__uuf__._1502_/X __dut__._2267_/B
+ __dut__.__uuf__._1491_/X __dut__.__uuf__._1509_/X VGND VGND VPWR VPWR __dut__._2266_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_116_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1441_ __dut__.__uuf__._1441_/A VGND VGND VPWR VPWR __dut__.__uuf__._1563_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1372_ __dut__._2327_/B VGND VGND VPWR VPWR __dut__.__uuf__._1372_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_143_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1692__A2 prod[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1444__A2 mc[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2040_ __dut__._2044_/A1 prod[2] __dut__._2039_/X VGND VGND VPWR VPWR __dut__._3077_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_26_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1264__B1 __dut__._2239_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1708_ __dut__.__uuf__._1699_/A __dut__.__uuf__._1706_/B __dut__.__uuf__._1661_/X
+ VGND VGND VPWR VPWR __dut__._2130_/A2 sky130_fd_sc_hd__o21a_4
X__dut__._2942_ __dut__._2958_/CLK __dut__._2942_/D __dut__._2676_/Y VGND VGND VPWR
+ VPWR __dut__._2942_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1639_ __dut__.__uuf__._1639_/A VGND VGND VPWR VPWR __dut__.__uuf__._1639_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2873_ clkbuf_5_9_0_tck/X __dut__._2873_/D __dut__._2745_/Y VGND VGND VPWR
+ VPWR __dut__._2873_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1031__A3 prod[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1824_ __dut__._1830_/A1 tie[64] __dut__._1823_/X VGND VGND VPWR VPWR __dut__._2969_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1380__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1755_ __dut__._2189_/A __dut__._2934_/Q VGND VGND VPWR VPWR __dut__._1755_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_150_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1686_ __dut__._1686_/A1 prod[60] __dut__._1685_/X VGND VGND VPWR VPWR __dut__._2900_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2307_ __dut__._2325_/A __dut__._2307_/B VGND VGND VPWR VPWR __dut__._2307_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2238_ __dut__._2238_/A1 __dut__._2238_/A2 __dut__._2237_/X VGND VGND VPWR
+ VPWR __dut__._2238_/X sky130_fd_sc_hd__a21o_4
X__dut__._2169_ __dut__._2207_/A __dut__._2169_/B VGND VGND VPWR VPWR __dut__._2169_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_240_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1990_ __dut__.__uuf__._1990_/A VGND VGND VPWR VPWR __dut__.__uuf__._1990_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_63_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1424_ __dut__.__uuf__._1422_/Y __dut__.__uuf__._1423_/X __dut__.__uuf__._1322_/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._1424_/X sky130_fd_sc_hd__o21a_4
XFILLER_144_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1355_ __dut__.__uuf__._1352_/X __dut__.__uuf__._1354_/X __dut__._2333_/B
+ __dut__.__uuf__._1352_/X VGND VGND VPWR VPWR __dut__._2332_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1540_ __dut__._1374_/Y mp[15] __dut__._1539_/X VGND VGND VPWR VPWR __dut__._1540_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1286_ __dut__.__uuf__._1308_/A VGND VGND VPWR VPWR __dut__.__uuf__._1286_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1471_ __dut__._2509_/A __dut__._2834_/Q VGND VGND VPWR VPWR __dut__._1471_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3072_ clkbuf_5_5_0_tck/X __dut__._3072_/D __dut__._2546_/Y VGND VGND VPWR
+ VPWR __dut__._3072_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1403__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2023_ __dut__._2207_/A __dut__._3068_/Q VGND VGND VPWR VPWR __dut__._2023_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_281_ _313_/CLK _281_/D VGND VGND VPWR VPWR _281_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__.__uuf__._1035__A __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_24_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2925_ clkbuf_5_9_0_tck/X __dut__._2925_/D __dut__._2693_/Y VGND VGND VPWR
+ VPWR __dut__._2925_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2856_ __dut__._2860_/CLK __dut__._2856_/D __dut__._2762_/Y VGND VGND VPWR
+ VPWR __dut__._2856_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1807_ __dut__._1807_/A __dut__._2960_/Q VGND VGND VPWR VPWR __dut__._1807_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2269__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2787_ rst VGND VGND VPWR VPWR __dut__._2787_/Y sky130_fd_sc_hd__inv_2
X__dut__._1738_ __dut__._1760_/A1 tie[21] __dut__._1737_/X VGND VGND VPWR VPWR __dut__._2926_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1669_ __dut__._2491_/A __dut__._2891_/Q VGND VGND VPWR VPWR __dut__._1669_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1408__A2 mc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1592__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_288_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1983__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1140_ __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR __dut__.__uuf__._1200_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1071_ __dut__.__uuf__._1071_/A VGND VGND VPWR VPWR __dut__.__uuf__._1071_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2319__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1973_ __dut__.__uuf__._1973_/A VGND VGND VPWR VPWR __dut__.__uuf__._1975_/B
+ sky130_fd_sc_hd__inv_2
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2710_ rst VGND VGND VPWR VPWR __dut__._2710_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1893__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2641_ rst VGND VGND VPWR VPWR __dut__._2641_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1407_ __dut__.__uuf__._1411_/A VGND VGND VPWR VPWR __dut__.__uuf__._1407_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_116_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2572_ rst VGND VGND VPWR VPWR __dut__._2572_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1338_ __dut__.__uuf__._1378_/A VGND VGND VPWR VPWR __dut__.__uuf__._1338_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2501__B prod[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1523_ __dut__._2509_/A __dut__._2847_/Q VGND VGND VPWR VPWR __dut__._1523_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1638__A2 prod[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1269_ __dut__.__uuf__._1266_/Y __dut__.__uuf__._1988_/B __dut__.__uuf__._1268_/X
+ VGND VGND VPWR VPWR __dut__._2364_/A2 sky130_fd_sc_hd__o21ai_4
XFILLER_100_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1454_ __dut__._2222_/A1 __dut__._1452_/X __dut__._1453_/X VGND VGND VPWR
+ VPWR __dut__._2829_/D sky130_fd_sc_hd__a21o_4
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1385_ __dut__._2189_/A __dut__._2811_/Q VGND VGND VPWR VPWR __dut__._1385_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2229__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._3055_ __dut__._3059_/CLK __dut__._3055_/D __dut__._2563_/Y VGND VGND VPWR
+ VPWR __dut__._3055_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2006_ __dut__._2006_/A1 tie[155] __dut__._2005_/X VGND VGND VPWR VPWR __dut__._3060_/D
+ sky130_fd_sc_hd__a21o_4
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_264_ _194_/A _264_/D VGND VGND VPWR VPWR _264_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_195_ _203_/A VGND VGND VPWR VPWR _199_/A sky130_fd_sc_hd__buf_2
XFILLER_127_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2908_ clkbuf_5_2_0_tck/X __dut__._2908_/D __dut__._2710_/Y VGND VGND VPWR
+ VPWR __dut__._2908_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_142_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2839_ __dut__._2846_/CLK __dut__._2839_/D __dut__._2779_/Y VGND VGND VPWR
+ VPWR __dut__._2839_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2054__A2 prod[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_203_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_14_0_tck clkbuf_4_7_0_tck/X VGND VGND VPWR VPWR __dut__._2958_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2310_ __dut__.__uuf__._2334_/CLK __dut__._2400_/X __dut__.__uuf__._1187_/X
+ VGND VGND VPWR VPWR prod[9] sky130_fd_sc_hd__dfrtp_4
XFILLER_127_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2241_ __dut__.__uuf__._2251_/CLK __dut__._2262_/X __dut__.__uuf__._1516_/X
+ VGND VGND VPWR VPWR __dut__._2263_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2602__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__312__SET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_29_0_tck clkbuf_5_29_0_tck/A VGND VGND VPWR VPWR __dut__._3059_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2172_ __dut__.__uuf__._2278_/CLK __dut__._2124_/X __dut__.__uuf__._1636_/X
+ VGND VGND VPWR VPWR __dut__._2125_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1123_ __dut__.__uuf__._1131_/A VGND VGND VPWR VPWR __dut__.__uuf__._1123_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1054_ __dut__.__uuf__._1099_/A VGND VGND VPWR VPWR __dut__.__uuf__._1054_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_56_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2049__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1956_ __dut__.__uuf__._1956_/A VGND VGND VPWR VPWR __dut__._2224_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_1_1_0_tck_A clkbuf_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1887_ __dut__._2199_/B __dut__._2205_/B __dut__.__uuf__._1886_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1888_/C sky130_fd_sc_hd__o21ai_4
XFILLER_137_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1556__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2821__CLK __dut__._2860_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2512__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2624_ rst VGND VGND VPWR VPWR __dut__._2624_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2555_ rst VGND VGND VPWR VPWR __dut__._2555_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_91_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1506_ __dut__._1506_/A1 __dut__._1504_/X __dut__._1505_/X VGND VGND VPWR
+ VPWR __dut__._2842_/D sky130_fd_sc_hd__a21o_4
XFILLER_143_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2486_ __dut__._2488_/A1 __dut__._2486_/A2 __dut__._2485_/X VGND VGND VPWR
+ VPWR __dut__._2486_/X sky130_fd_sc_hd__a21o_4
X__dut__._1437_ __dut__._1437_/A __dut__._2824_/Q VGND VGND VPWR VPWR __dut__._1437_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._3107_ __dut__._3109_/CLK __dut__._3107_/D __dut__._2511_/Y VGND VGND VPWR
+ VPWR __dut__._3107_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3038_ _306_/CLK __dut__._3038_/D __dut__._2580_/Y VGND VGND VPWR VPWR __dut__._3038_/Q
+ sky130_fd_sc_hd__dfrtp_4
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_247_ _202_/X _311_/Q VGND VGND VPWR VPWR _247_/Q sky130_fd_sc_hd__dfxtp_4
X_178_ _274_/Q _182_/B VGND VGND VPWR VPWR _273_/D sky130_fd_sc_hd__and2_4
XFILLER_143_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_153_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1810_ __dut__._2171_/B __dut__._2177_/B __dut__.__uuf__._1809_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1811_/C sky130_fd_sc_hd__o21ai_4
XANTENNA__268__CLK _274_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1741_ __dut__.__uuf__._1734_/A __dut__.__uuf__._1739_/B __dut__.__uuf__._1720_/X
+ VGND VGND VPWR VPWR __dut__._2142_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_119_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1672_ __dut__.__uuf__._1261_/X __dut__.__uuf__._1670_/B __dut__.__uuf__._1670_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1673_/C sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._1501__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2844__CLK __dut__._2846_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2994__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2224_ __dut__.__uuf__._2291_/CLK __dut__._2228_/X __dut__.__uuf__._1571_/X
+ VGND VGND VPWR VPWR __dut__._2229_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2155_ VGND VGND VPWR VPWR __dut__.__uuf__._2155_/HI tie[162] sky130_fd_sc_hd__conb_1
XFILLER_102_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1106_ __dut__.__uuf__._1117_/A VGND VGND VPWR VPWR __dut__.__uuf__._1106_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_113_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2340_ __dut__._2368_/A1 __dut__._2340_/A2 __dut__._2339_/X VGND VGND VPWR
+ VPWR __dut__._2340_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2086_ VGND VGND VPWR VPWR __dut__.__uuf__._2086_/HI tie[93] sky130_fd_sc_hd__conb_1
X__dut__._2271_ __dut__._2281_/A __dut__._2271_/B VGND VGND VPWR VPWR __dut__._2271_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1037_ __dut__.__uuf__._1019_/X __dut__.__uuf__._1023_/X prod[60]
+ prod[61] __dut__.__uuf__._1036_/X VGND VGND VPWR VPWR __dut__._2502_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1939_ __dut__._2219_/B __dut__._2225_/B VGND VGND VPWR VPWR __dut__.__uuf__._1940_/A
+ sky130_fd_sc_hd__and2_4
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2507__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1411__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1986_ __dut__._2004_/A1 tie[145] __dut__._1985_/X VGND VGND VPWR VPWR __dut__._3050_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_152_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2607_ rst VGND VGND VPWR VPWR __dut__._2607_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2538_ rst VGND VGND VPWR VPWR __dut__._2538_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2469_ __dut__._2491_/A prod[43] VGND VGND VPWR VPWR __dut__._2469_/X sky130_fd_sc_hd__and2_4
XFILLER_74_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_270_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1991__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2327__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1724_ __dut__.__uuf__._1724_/A VGND VGND VPWR VPWR __dut__.__uuf__._1724_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_33_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._3022__CLK clkbuf_opt_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1655_ __dut__._2111_/B __dut__._2121_/B __dut__.__uuf__._1654_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1656_/C sky130_fd_sc_hd__o21ai_4
XFILLER_147_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1840_ __dut__._1840_/A1 tie[72] __dut__._1839_/X VGND VGND VPWR VPWR __dut__._2977_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1586_ __dut__.__uuf__._1590_/A VGND VGND VPWR VPWR __dut__.__uuf__._1586_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_108_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1771_ __dut__._1775_/A __dut__._2942_/Q VGND VGND VPWR VPWR __dut__._1771_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2207_ __dut__.__uuf__._2230_/CLK __dut__._2194_/X __dut__.__uuf__._1593_/X
+ VGND VGND VPWR VPWR __dut__._2195_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_76_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2138_ VGND VGND VPWR VPWR __dut__.__uuf__._2138_/HI tie[145] sky130_fd_sc_hd__conb_1
XFILLER_124_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__245__A1 tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2323_ __dut__._2325_/A __dut__._2323_/B VGND VGND VPWR VPWR __dut__._2323_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._2069_ VGND VGND VPWR VPWR __dut__.__uuf__._2069_/HI tie[76] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._1998__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2254_ __dut__._2256_/A1 __dut__._2254_/A2 __dut__._2253_/X VGND VGND VPWR
+ VPWR __dut__._2254_/X sky130_fd_sc_hd__a21o_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_103 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1786_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2185_ __dut__._2189_/A __dut__._2185_/B VGND VGND VPWR VPWR __dut__._2185_/X
+ sky130_fd_sc_hd__and2_4
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_4_0_tck clkbuf_4_5_0_tck/A VGND VGND VPWR VPWR clkbuf_5_9_0_tck/A sky130_fd_sc_hd__clkbuf_1
Xpsn_inst_psn_buff_136 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2074_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_114 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1836_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_125 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1870_/A1 sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2237__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_147 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2440_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_158 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2450_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_169 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2004_/A1 sky130_fd_sc_hd__buf_8
XFILLER_149_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1969_ __dut__._1969_/A __dut__._3041_/Q VGND VGND VPWR VPWR __dut__._1969_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_4_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2700__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._3045__CLK __dut__._3058_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_116_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2147__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1440_ __dut__.__uuf__._1463_/A VGND VGND VPWR VPWR __dut__.__uuf__._1440_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2166__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1371_ __dut__.__uuf__._1386_/A VGND VGND VPWR VPWR __dut__.__uuf__._1371_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_104_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_0_0_tck_A clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2610__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_7_0___dut__.__uuf__.__clk_source__ clkbuf_4_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2278_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1264__B2 __dut__.__uuf__._1025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2057__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1707_ __dut__.__uuf__._1707_/A VGND VGND VPWR VPWR __dut__._2132_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__._2941_ __dut__._2941_/CLK __dut__._2941_/D __dut__._2677_/Y VGND VGND VPWR
+ VPWR __dut__._2941_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1638_ __dut__.__uuf__._1639_/A VGND VGND VPWR VPWR __dut__.__uuf__._1638_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1904__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2872_ clkbuf_5_2_0_tck/X __dut__._2872_/D __dut__._2746_/Y VGND VGND VPWR
+ VPWR __dut__._2872_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1823_ __dut__._2507_/A __dut__._2968_/Q VGND VGND VPWR VPWR __dut__._1823_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1569_ __dut__.__uuf__._1571_/A VGND VGND VPWR VPWR __dut__.__uuf__._1569_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1754_ __dut__._1760_/A1 tie[29] __dut__._1753_/X VGND VGND VPWR VPWR __dut__._2934_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1380__A2 mc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2520__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1685_ __dut__._2503_/A __dut__._2899_/Q VGND VGND VPWR VPWR __dut__._1685_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_135_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._3068__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2306_ __dut__._2308_/A1 __dut__._2306_/A2 __dut__._2305_/X VGND VGND VPWR
+ VPWR __dut__._2306_/X sky130_fd_sc_hd__a21o_4
X__dut__._2237_ __dut__._2325_/A __dut__._2237_/B VGND VGND VPWR VPWR __dut__._2237_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2198__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2168_ __dut__._2172_/A1 __dut__._2168_/A2 __dut__._2167_/X VGND VGND VPWR
+ VPWR __dut__._2168_/X sky130_fd_sc_hd__a21o_4
XFILLER_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2396__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2099_ __dut__._2507_/A __dut__._3106_/Q VGND VGND VPWR VPWR __dut__._2099_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2320__A1 __dut__._2332_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_233_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2605__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1423_ __dut__.__uuf__._1492_/A VGND VGND VPWR VPWR __dut__.__uuf__._1423_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_144_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1354_ __dut__.__uuf__._1353_/Y __dut__.__uuf__._1347_/X __dut__.__uuf__._1348_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1354_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1285_ __dut__.__uuf__._1340_/A VGND VGND VPWR VPWR __dut__.__uuf__._1308_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_98_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1470_ __dut__._1474_/A1 __dut__._1468_/X __dut__._1469_/X VGND VGND VPWR
+ VPWR __dut__._2833_/D sky130_fd_sc_hd__a21o_4
XFILLER_86_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3071_ clkbuf_5_5_0_tck/X __dut__._3071_/D __dut__._2547_/Y VGND VGND VPWR
+ VPWR __dut__._3071_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2022_ __dut__._2022_/A1 tie[163] __dut__._2021_/X VGND VGND VPWR VPWR __dut__._3068_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_280_ _194_/A _280_/D VGND VGND VPWR VPWR _280_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._2378__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_17_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2515__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2924_ clkbuf_5_9_0_tck/X __dut__._2924_/D __dut__._2694_/Y VGND VGND VPWR
+ VPWR __dut__._2924_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1051__A __dut__.__uuf__._1214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2855_ __dut__._2860_/CLK __dut__._2855_/D __dut__._2763_/Y VGND VGND VPWR
+ VPWR __dut__._2855_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1806_ __dut__._1806_/A1 tie[55] __dut__._1805_/X VGND VGND VPWR VPWR __dut__._2960_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2786_ rst VGND VGND VPWR VPWR __dut__._2786_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1737_ __dut__._2189_/A __dut__._2925_/Q VGND VGND VPWR VPWR __dut__._1737_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1668_ __dut__._2488_/A1 prod[51] __dut__._1667_/X VGND VGND VPWR VPWR __dut__._2891_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1599_ __dut__._2509_/A __dut__._2866_/Q VGND VGND VPWR VPWR __dut__._1599_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_91_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2425__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1592__A2 mp[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2213__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_113_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1070_ __dut__.__uuf__._1057_/X __dut__.__uuf__._1069_/X prod[49]
+ prod[50] __dut__.__uuf__._1066_/X VGND VGND VPWR VPWR __dut__._2480_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_95_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1972_ __dut__.__uuf__._1982_/A __dut__.__uuf__._1972_/B __dut__.__uuf__._1972_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1973_/A sky130_fd_sc_hd__or3_4
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2335__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2640_ rst VGND VGND VPWR VPWR __dut__._2640_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1406_ __dut__.__uuf__._1403_/X __dut__.__uuf__._1405_/X __dut__._2313_/B
+ __dut__.__uuf__._1403_/X VGND VGND VPWR VPWR __dut__._2312_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1337_ __dut__.__uuf__._1336_/Y __dut__.__uuf__._1321_/X __dut__.__uuf__._1322_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1337_/X sky130_fd_sc_hd__o21a_4
X__dut__._2571_ rst VGND VGND VPWR VPWR __dut__._2571_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1522_ __dut__._1522_/A1 __dut__._1520_/X __dut__._1521_/X VGND VGND VPWR
+ VPWR __dut__._2846_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1268_ __dut__.__uuf__._1399_/A VGND VGND VPWR VPWR __dut__.__uuf__._1268_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_74_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1199_ __dut__.__uuf__._1205_/A VGND VGND VPWR VPWR __dut__.__uuf__._1199_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1453_ __dut__._2325_/A __dut__._2828_/Q VGND VGND VPWR VPWR __dut__._1453_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_132_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1384_ __dut__._1374_/Y mc[11] __dut__._1383_/X VGND VGND VPWR VPWR __dut__._1384_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_54_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._3054_ __dut__._3059_/CLK __dut__._3054_/D __dut__._2564_/Y VGND VGND VPWR
+ VPWR __dut__._3054_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._3106__CLK __dut__._3106_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2005_ __dut__._2005_/A __dut__._3059_/Q VGND VGND VPWR VPWR __dut__._2005_/X
+ sky130_fd_sc_hd__and2_4
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_263_ _194_/A _263_/D VGND VGND VPWR VPWR _263_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_194_ _194_/A VGND VGND VPWR VPWR _203_/A sky130_fd_sc_hd__inv_2
XFILLER_6_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2236__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2907_ clkbuf_5_2_0_tck/X __dut__._2907_/D __dut__._2711_/Y VGND VGND VPWR
+ VPWR __dut__._2907_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2838_ __dut__._2846_/CLK __dut__._2838_/D __dut__._2780_/Y VGND VGND VPWR
+ VPWR __dut__._2838_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2769_ rst VGND VGND VPWR VPWR __dut__._2769_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2155__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2240_ __dut__.__uuf__._2240_/CLK __dut__._2260_/X __dut__.__uuf__._1519_/X
+ VGND VGND VPWR VPWR __dut__._2261_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2171_ __dut__.__uuf__._2278_/CLK __dut__._2122_/X __dut__.__uuf__._1637_/X
+ VGND VGND VPWR VPWR __dut__._2123_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1122_ __dut__.__uuf__._1118_/X __dut__.__uuf__._1115_/X prod[32]
+ prod[33] __dut__.__uuf__._1111_/X VGND VGND VPWR VPWR __dut__._2446_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_101_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_10_0_tck_A clkbuf_3_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1053_ __dut__.__uuf__._1056_/A VGND VGND VPWR VPWR __dut__.__uuf__._1053_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1955_ __dut__.__uuf__._1975_/A __dut__.__uuf__._1955_/B __dut__.__uuf__._1955_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1956_/A sky130_fd_sc_hd__or3_4
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1886_ __dut__.__uuf__._1886_/A VGND VGND VPWR VPWR __dut__.__uuf__._1886_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_137_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1556__A2 mp[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__213__A tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1409__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2623_ rst VGND VGND VPWR VPWR __dut__._2623_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2554_ rst VGND VGND VPWR VPWR __dut__._2554_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_84_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1505_ __dut__._2189_/A __dut__._2841_/Q VGND VGND VPWR VPWR __dut__._1505_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_143_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2485_ __dut__._2491_/A prod[51] VGND VGND VPWR VPWR __dut__._2485_/X sky130_fd_sc_hd__and2_4
XFILLER_74_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1492__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1436_ __dut__._1374_/Y mc[23] __dut__._1435_/X VGND VGND VPWR VPWR __dut__._1436_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._3106_ __dut__._3106_/CLK __dut__._3106_/D __dut__._2512_/Y VGND VGND VPWR
+ VPWR __dut__._3106_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3037_ _290_/CLK __dut__._3037_/D __dut__._2581_/Y VGND VGND VPWR VPWR __dut__._3037_/Q
+ sky130_fd_sc_hd__dfrtp_4
X_315_ _315_/CLK _315_/D trst VGND VGND VPWR VPWR _315_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_246_ _203_/X _295_/Q VGND VGND VPWR VPWR _246_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_177_ _275_/Q _182_/B VGND VGND VPWR VPWR _274_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2703__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1119__B1 prod[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_146_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1989__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._1740_ __dut__.__uuf__._1740_/A VGND VGND VPWR VPWR __dut__._2144_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_119_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1671_ __dut__.__uuf__._1671_/A VGND VGND VPWR VPWR __dut__.__uuf__._1673_/B
+ sky130_fd_sc_hd__inv_2
Xclkbuf_3_0_0___dut__.__uuf__.__clk_source__ clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_1_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_107_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2613__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2223_ __dut__.__uuf__._2225_/CLK __dut__._2226_/X __dut__.__uuf__._1574_/X
+ VGND VGND VPWR VPWR __dut__._2227_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_142_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2154_ VGND VGND VPWR VPWR __dut__.__uuf__._2154_/HI tie[161] sky130_fd_sc_hd__conb_1
XFILLER_102_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1105_ __dut__.__uuf__._1134_/A VGND VGND VPWR VPWR __dut__.__uuf__._1117_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2085_ VGND VGND VPWR VPWR __dut__.__uuf__._2085_/HI tie[92] sky130_fd_sc_hd__conb_1
XFILLER_113_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2270_ __dut__._2278_/A1 __dut__._2270_/A2 __dut__._2269_/X VGND VGND VPWR
+ VPWR __dut__._2270_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1036_ __dut__.__uuf__._1214_/A VGND VGND VPWR VPWR __dut__.__uuf__._1036_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1899__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1938_ __dut__._1448_/X VGND VGND VPWR VPWR __dut__.__uuf__._1942_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2507__B prod[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1869_ __dut__.__uuf__._1869_/A __dut__.__uuf__._1869_/B __dut__.__uuf__._1869_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1870_/A sky130_fd_sc_hd__or3_4
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1985_ __dut__._2005_/A __dut__._3049_/Q VGND VGND VPWR VPWR __dut__._1985_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2523__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2606_ rst VGND VGND VPWR VPWR __dut__._2606_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1116__A3 prod[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2537_ rst VGND VGND VPWR VPWR __dut__._2537_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2468_ __dut__._2488_/A1 __dut__._2468_/A2 __dut__._2467_/X VGND VGND VPWR
+ VPWR __dut__._2468_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_13_0_tck clkbuf_4_6_0_tck/X VGND VGND VPWR VPWR __dut__._2860_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__._1419_ __dut__._2509_/A __dut__._2821_/Q VGND VGND VPWR VPWR __dut__._1419_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_35_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2399_ __dut__._2407_/A prod[8] VGND VGND VPWR VPWR __dut__._2399_/X sky130_fd_sc_hd__and2_4
XFILLER_97_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_28_0_tck clkbuf_5_29_0_tck/A VGND VGND VPWR VPWR _271_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_229_ _299_/Q _228_/B _222_/A VGND VGND VPWR VPWR _302_/D sky130_fd_sc_hd__o21a_4
XFILLER_144_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2433__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_263_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1107__A3 prod[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1456__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2608__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1723_ __dut__._2139_/B __dut__._2145_/B VGND VGND VPWR VPWR __dut__.__uuf__._1724_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_138_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1654_ __dut__.__uuf__._1654_/A VGND VGND VPWR VPWR __dut__.__uuf__._1654_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_119_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1585_ __dut__.__uuf__._1597_/A VGND VGND VPWR VPWR __dut__.__uuf__._1590_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2343__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1770_ __dut__._1780_/A1 tie[37] __dut__._1769_/X VGND VGND VPWR VPWR __dut__._2942_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_108_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2206_ __dut__.__uuf__._2230_/CLK __dut__._2192_/X __dut__.__uuf__._1594_/X
+ VGND VGND VPWR VPWR __dut__._2193_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_124_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2137_ VGND VGND VPWR VPWR __dut__.__uuf__._2137_/HI tie[144] sky130_fd_sc_hd__conb_1
XFILLER_124_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2322_ __dut__._2332_/A1 __dut__._2322_/A2 __dut__._2321_/X VGND VGND VPWR
+ VPWR __dut__._2322_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2068_ VGND VGND VPWR VPWR __dut__.__uuf__._2068_/HI tie[75] sky130_fd_sc_hd__conb_1
XFILLER_72_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1019_ __dut__.__uuf__._1088_/A VGND VGND VPWR VPWR __dut__.__uuf__._1019_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_140_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2253_ __dut__._2253_/A __dut__._2253_/B VGND VGND VPWR VPWR __dut__._2253_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2518__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2184_ __dut__._2184_/A1 __dut__._2184_/A2 __dut__._2183_/X VGND VGND VPWR
+ VPWR __dut__._2184_/X sky130_fd_sc_hd__a21o_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_137 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2424_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_104 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1788_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_126 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1872_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_115 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1838_/A1 sky130_fd_sc_hd__buf_2
XFILLER_25_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_148 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2094_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_159 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2104_/A1 sky130_fd_sc_hd__buf_2
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1968_ __dut__._2004_/A1 tie[136] __dut__._1967_/X VGND VGND VPWR VPWR __dut__._3041_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_140_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1899_ __dut__._2005_/A __dut__._3006_/Q VGND VGND VPWR VPWR __dut__._1899_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1229__A __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_109_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__301__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2163__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1370_ __dut__.__uuf__._1363_/X __dut__.__uuf__._1369_/X __dut__._2327_/B
+ __dut__.__uuf__._1363_/X VGND VGND VPWR VPWR __dut__._2326_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1507__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1706_ __dut__.__uuf__._1706_/A __dut__.__uuf__._1706_/B __dut__.__uuf__._1706_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1707_/A sky130_fd_sc_hd__or3_4
X__dut__._2940_ __dut__._2941_/CLK __dut__._2940_/D __dut__._2678_/Y VGND VGND VPWR
+ VPWR __dut__._2940_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1637_ __dut__.__uuf__._1639_/A VGND VGND VPWR VPWR __dut__.__uuf__._1637_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2871_ clkbuf_5_3_0_tck/X __dut__._2871_/D __dut__._2747_/Y VGND VGND VPWR
+ VPWR __dut__._2871_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1822_ __dut__._1830_/A1 tie[63] __dut__._1821_/X VGND VGND VPWR VPWR __dut__._2968_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1568_ __dut__.__uuf__._1571_/A VGND VGND VPWR VPWR __dut__.__uuf__._1568_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1753_ __dut__._2189_/A __dut__._2933_/Q VGND VGND VPWR VPWR __dut__._1753_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2801__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1499_ __dut__._1544_/X __dut__.__uuf__._1487_/X __dut__._2273_/B
+ __dut__.__uuf__._1492_/X VGND VGND VPWR VPWR __dut__.__uuf__._1499_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__._2857__CLK __dut__._2860_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1668__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1684_ __dut__._2004_/A1 prod[59] __dut__._1683_/X VGND VGND VPWR VPWR __dut__._2899_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_135_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1417__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2305_ __dut__._2325_/A __dut__._2305_/B VGND VGND VPWR VPWR __dut__._2305_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2236_ __dut__._2236_/A1 __dut__._2236_/A2 __dut__._2235_/X VGND VGND VPWR
+ VPWR __dut__._2236_/X sky130_fd_sc_hd__a21o_4
XFILLER_32_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2167_ __dut__._2207_/A __dut__._2167_/B VGND VGND VPWR VPWR __dut__._2167_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2098_ __dut__._2098_/A1 prod[31] __dut__._2097_/X VGND VGND VPWR VPWR __dut__._3106_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_138_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1512__A __dut__.__uuf__._1533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2711__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3012__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2084__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_226_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1997__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1422_ __dut__._2307_/B VGND VGND VPWR VPWR __dut__.__uuf__._1422_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_116_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1898__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1353_ __dut__._2335_/B VGND VGND VPWR VPWR __dut__.__uuf__._1353_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2621__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_3_0_tck clkbuf_4_3_0_tck/A VGND VGND VPWR VPWR clkbuf_5_7_0_tck/A sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1284_ __dut__.__uuf__._1271_/X __dut__.__uuf__._1282_/X __dut__._2359_/B
+ __dut__.__uuf__._1283_/X VGND VGND VPWR VPWR __dut__._2358_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3070_ clkbuf_5_5_0_tck/X __dut__._3070_/D __dut__._2548_/Y VGND VGND VPWR
+ VPWR __dut__._3070_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2021_ __dut__._2207_/A __dut__._3067_/Q VGND VGND VPWR VPWR __dut__._2021_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__294__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2923_ clkbuf_5_9_0_tck/X __dut__._2923_/D __dut__._2695_/Y VGND VGND VPWR
+ VPWR __dut__._2923_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2854_ clkbuf_5_3_0_tck/X __dut__._2854_/D __dut__._2764_/Y VGND VGND VPWR
+ VPWR __dut__._2854_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1805_ __dut__._1805_/A __dut__._2959_/Q VGND VGND VPWR VPWR __dut__._1805_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2785_ rst VGND VGND VPWR VPWR __dut__._2785_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2531__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3035__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1736_ __dut__._1760_/A1 tie[20] __dut__._1735_/X VGND VGND VPWR VPWR __dut__._2925_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1667_ __dut__._2491_/A __dut__._2890_/Q VGND VGND VPWR VPWR __dut__._1667_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_130_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1598_ __dut__._1598_/A1 __dut__._1596_/X __dut__._1597_/X VGND VGND VPWR
+ VPWR __dut__._2865_/D sky130_fd_sc_hd__a21o_4
XFILLER_76_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2066__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2165__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_91_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1507__A __dut__.__uuf__._1549_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2219_ __dut__._2325_/A __dut__._2219_/B VGND VGND VPWR VPWR __dut__._2219_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2706__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2441__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_176_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1971_ __dut__._2231_/B __dut__._2237_/B __dut__.__uuf__._1970_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1972_/C sky130_fd_sc_hd__o21ai_4
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2616__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3058__CLK __dut__._3058_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2351__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1405_ __dut__.__uuf__._1404_/Y __dut__.__uuf__._1398_/X __dut__.__uuf__._1399_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1405_/X sky130_fd_sc_hd__o21a_4
XFILLER_105_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1336_ __dut__._2341_/B VGND VGND VPWR VPWR __dut__.__uuf__._1336_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._2570_ rst VGND VGND VPWR VPWR __dut__._2570_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__.__uuf__._2188__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1521_ __dut__._1557_/A __dut__._2845_/Q VGND VGND VPWR VPWR __dut__._1521_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1267_ __dut__._1612_/X __dut__.__uuf__._1292_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1399_/A sky130_fd_sc_hd__nand2_4
XFILLER_112_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1198_ __dut__.__uuf__._1192_/X __dut__.__uuf__._1189_/X prod[6]
+ prod[7] __dut__.__uuf__._1185_/X VGND VGND VPWR VPWR __dut__._2394_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1452_ __dut__._1374_/Y mc[27] __dut__._1451_/X VGND VGND VPWR VPWR __dut__._1452_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_132_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1383_ __dut__._2509_/A __dut__._2812_/Q VGND VGND VPWR VPWR __dut__._1383_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2048__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3053_ __dut__._3059_/CLK __dut__._3053_/D __dut__._2565_/Y VGND VGND VPWR
+ VPWR __dut__._3053_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2004_ __dut__._2004_/A1 tie[154] __dut__._2003_/X VGND VGND VPWR VPWR __dut__._3059_/D
+ sky130_fd_sc_hd__a21o_4
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2526__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_262_ _194_/A _262_/D VGND VGND VPWR VPWR _262_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_193_ _260_/Q _193_/B VGND VGND VPWR VPWR _259_/D sky130_fd_sc_hd__or2_4
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._2906_ clkbuf_5_0_0_tck/X __dut__._2906_/D __dut__._2712_/Y VGND VGND VPWR
+ VPWR __dut__._2906_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2837_ __dut__._2846_/CLK __dut__._2837_/D __dut__._2781_/Y VGND VGND VPWR
+ VPWR __dut__._2837_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2768_ rst VGND VGND VPWR VPWR __dut__._2768_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1719_ __dut__._2189_/A __dut__._2916_/Q VGND VGND VPWR VPWR __dut__._1719_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2699_ rst VGND VGND VPWR VPWR __dut__._2699_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1237__A __dut__.__uuf__._1640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1970__B1 __dut__._1969_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_293_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2171__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2170_ __dut__.__uuf__._2278_/CLK __dut__._2120_/X __dut__.__uuf__._1638_/X
+ VGND VGND VPWR VPWR __dut__._2121_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_142_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1121_ __dut__.__uuf__._1131_/A VGND VGND VPWR VPWR __dut__.__uuf__._1121_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_68_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1052_ __dut__.__uuf__._1043_/X __dut__.__uuf__._1040_/X prod[55]
+ prod[56] __dut__.__uuf__._1051_/X VGND VGND VPWR VPWR __dut__._2492_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1515__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1954_ __dut__.__uuf__._1921_/X __dut__.__uuf__._1952_/B __dut__.__uuf__._1952_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1955_/C sky130_fd_sc_hd__o21a_4
XFILLER_12_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1885_ __dut__._2199_/B __dut__._2205_/B VGND VGND VPWR VPWR __dut__.__uuf__._1886_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_137_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1610__A __dut__.__uuf__._1628_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2622_ rst VGND VGND VPWR VPWR __dut__._2622_/Y sky130_fd_sc_hd__inv_2
X__dut__._2553_ rst VGND VGND VPWR VPWR __dut__._2553_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2299_ __dut__.__uuf__._2303_/CLK __dut__._2378_/X __dut__.__uuf__._1234_/X
+ VGND VGND VPWR VPWR __dut__._2379_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1319_ __dut__._2347_/B VGND VGND VPWR VPWR __dut__.__uuf__._1319_/Y
+ sky130_fd_sc_hd__inv_2
Xclkbuf_opt_2_tck clkbuf_opt_2_tck/A VGND VGND VPWR VPWR clkbuf_opt_2_tck/X sky130_fd_sc_hd__clkbuf_16
X__dut__._1504_ __dut__._1374_/Y mp[7] __dut__._1503_/X VGND VGND VPWR VPWR __dut__._1504_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_101_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_77_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2484_ __dut__._2488_/A1 __dut__._2484_/A2 __dut__._2483_/X VGND VGND VPWR
+ VPWR __dut__._2484_/X sky130_fd_sc_hd__a21o_4
XFILLER_143_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1492__A2 mp[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1435_ __dut__._2509_/A __dut__._2825_/Q VGND VGND VPWR VPWR __dut__._1435_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3105_ __dut__._3106_/CLK __dut__._3105_/D __dut__._2513_/Y VGND VGND VPWR
+ VPWR __dut__._3105_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._3036_ clkbuf_5_4_0_tck/X __dut__._3036_/D __dut__._2582_/Y VGND VGND VPWR
+ VPWR __dut__._3036_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._2203__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_314_ _315_/CLK _314_/D trst VGND VGND VPWR VPWR _314_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_245_ tdi _154_/C _302_/Q _315_/Q VGND VGND VPWR VPWR _315_/D sky130_fd_sc_hd__o22a_4
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_176_ _183_/A VGND VGND VPWR VPWR _182_/B sky130_fd_sc_hd__buf_2
XFILLER_115_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_139_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1670_ __dut__.__uuf__._1680_/A __dut__.__uuf__._1670_/B __dut__.__uuf__._1670_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1671_/A sky130_fd_sc_hd__or3_4
XFILLER_146_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2222_ __dut__.__uuf__._2225_/CLK __dut__._2224_/X __dut__.__uuf__._1575_/X
+ VGND VGND VPWR VPWR __dut__._2225_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2153_ VGND VGND VPWR VPWR __dut__.__uuf__._2153_/HI tie[160] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2890__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1104_ __dut__.__uuf__._1103_/X __dut__.__uuf__._1099_/X prod[38]
+ prod[39] __dut__.__uuf__._1096_/X VGND VGND VPWR VPWR __dut__._2458_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2084_ VGND VGND VPWR VPWR __dut__.__uuf__._2084_/HI tie[91] sky130_fd_sc_hd__conb_1
XFILLER_113_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1035_ __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR __dut__.__uuf__._1214_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2226__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1937_ __dut__.__uuf__._1929_/A __dut__.__uuf__._1934_/B __dut__.__uuf__._1936_/X
+ VGND VGND VPWR VPWR __dut__._2214_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_138_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1868_ __dut__.__uuf__._1867_/X __dut__.__uuf__._1865_/B __dut__.__uuf__._1865_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1869_/C sky130_fd_sc_hd__o21a_4
XFILLER_149_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2804__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1934__B1 __dut__._1933_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1799_ __dut__.__uuf__._1799_/A VGND VGND VPWR VPWR __dut__.__uuf__._1799_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1984_ __dut__._2004_/A1 tie[144] __dut__._1983_/X VGND VGND VPWR VPWR __dut__._3049_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_106_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2605_ rst VGND VGND VPWR VPWR __dut__._2605_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2536_ rst VGND VGND VPWR VPWR __dut__._2536_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2467_ __dut__._2491_/A prod[42] VGND VGND VPWR VPWR __dut__._2467_/X sky130_fd_sc_hd__and2_4
X__dut__._1418_ __dut__._1418_/A1 __dut__._1416_/X __dut__._1417_/X VGND VGND VPWR
+ VPWR __dut__._2820_/D sky130_fd_sc_hd__a21o_4
X__dut__._2398_ __dut__._2412_/A1 __dut__._2398_/A2 __dut__._2397_/X VGND VGND VPWR
+ VPWR __dut__._2398_/X sky130_fd_sc_hd__a21o_4
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3019_ clkbuf_opt_2_tck/A __dut__._3019_/D __dut__._2599_/Y VGND VGND VPWR
+ VPWR __dut__._3019_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1037__B1 prod[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_228_ _232_/A _228_/B VGND VGND VPWR VPWR _301_/D sky130_fd_sc_hd__and2_4
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2714__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_159_ _289_/Q _164_/B VGND VGND VPWR VPWR _288_/D sky130_fd_sc_hd__and2_4
XFILLER_7_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_256_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1456__A2 mc[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1722_ __dut__._1620_/X VGND VGND VPWR VPWR __dut__.__uuf__._1726_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1653_ __dut__._2111_/B __dut__._2121_/B VGND VGND VPWR VPWR __dut__.__uuf__._1654_/A
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1916__B1 __dut__._1915_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2624__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1584_ __dut__.__uuf__._1584_/A VGND VGND VPWR VPWR __dut__.__uuf__._1584_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1392__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2205_ __dut__.__uuf__._2230_/CLK __dut__._2190_/X __dut__.__uuf__._1595_/X
+ VGND VGND VPWR VPWR __dut__._2191_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_103_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2136_ VGND VGND VPWR VPWR __dut__.__uuf__._2136_/HI tie[143] sky130_fd_sc_hd__conb_1
XFILLER_124_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2321_ __dut__._2325_/A __dut__._2321_/B VGND VGND VPWR VPWR __dut__._2321_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._2067_ VGND VGND VPWR VPWR __dut__.__uuf__._2067_/HI tie[74] sky130_fd_sc_hd__conb_1
X__dut__._2252_ __dut__._2256_/A1 __dut__._2252_/A2 __dut__._2251_/X VGND VGND VPWR
+ VPWR __dut__._2252_/X sky130_fd_sc_hd__a21o_4
XFILLER_17_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1018_ __dut__.__uuf__._1549_/A VGND VGND VPWR VPWR __dut__.__uuf__._1088_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1703__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2183_ __dut__._2189_/A __dut__._2183_/B VGND VGND VPWR VPWR __dut__._2183_/X
+ sky130_fd_sc_hd__and2_4
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_105 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1790_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_127 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1874_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_116 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1840_/A1 sky130_fd_sc_hd__buf_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_138 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2426_/A1 sky130_fd_sc_hd__buf_2
XFILLER_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_149 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2442_/A1 sky130_fd_sc_hd__buf_2
XFILLER_149_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__.__uuf__._1989__B __dut__._2109_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2534__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1967_ __dut__._1967_/A __dut__._3040_/Q VGND VGND VPWR VPWR __dut__._1967_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1898_ __dut__._2004_/A1 tie[101] __dut__._1897_/X VGND VGND VPWR VPWR __dut__._3006_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1686__A2 prod[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2519_ rst VGND VGND VPWR VPWR __dut__._2519_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2709__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3091__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1523__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2619__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1705_ __dut__.__uuf__._1704_/X __dut__.__uuf__._1701_/B __dut__.__uuf__._1701_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1706_/C sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1636_ __dut__.__uuf__._1639_/A VGND VGND VPWR VPWR __dut__.__uuf__._1636_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2870_ __dut__._2961_/CLK __dut__._2870_/D __dut__._2748_/Y VGND VGND VPWR
+ VPWR __dut__._2870_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1821_ __dut__._1821_/A __dut__._2967_/Q VGND VGND VPWR VPWR __dut__._1821_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1567_ __dut__.__uuf__._1571_/A VGND VGND VPWR VPWR __dut__.__uuf__._1567_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_123_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_12_0_tck clkbuf_4_6_0_tck/X VGND VGND VPWR VPWR __dut__._2941_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_134_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1752_ __dut__._1760_/A1 tie[28] __dut__._1751_/X VGND VGND VPWR VPWR __dut__._2933_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1498_ __dut__.__uuf__._1501_/A VGND VGND VPWR VPWR __dut__.__uuf__._1498_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1683_ __dut__._1891_/A __dut__._2898_/Q VGND VGND VPWR VPWR __dut__._1683_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_130_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_27_0_tck clkbuf_5_27_0_tck/A VGND VGND VPWR VPWR _194_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2119_ VGND VGND VPWR VPWR __dut__.__uuf__._2119_/HI tie[126] sky130_fd_sc_hd__conb_1
XFILLER_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2304_ __dut__._2308_/A1 __dut__._2304_/A2 __dut__._2303_/X VGND VGND VPWR
+ VPWR __dut__._2304_/X sky130_fd_sc_hd__a21o_4
XFILLER_57_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1433__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2529__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2235_ __dut__._2325_/A __dut__._2235_/B VGND VGND VPWR VPWR __dut__._2235_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_44_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1065__A __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2166_ __dut__._2172_/A1 __dut__._2166_/A2 __dut__._2165_/X VGND VGND VPWR
+ VPWR __dut__._2166_/X sky130_fd_sc_hd__a21o_4
X__dut__._2097_ __dut__._2507_/A __dut__._3105_/Q VGND VGND VPWR VPWR __dut__._2097_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2999_ __dut__._3096_/CLK __dut__._2999_/D __dut__._2619_/Y VGND VGND VPWR
+ VPWR __dut__._2999_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2439__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_121_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_219_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1421_ __dut__.__uuf__._1434_/A VGND VGND VPWR VPWR __dut__.__uuf__._1421_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_116_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1352_ __dut__.__uuf__._1378_/A VGND VGND VPWR VPWR __dut__.__uuf__._1352_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1283_ __dut__.__uuf__._1311_/A VGND VGND VPWR VPWR __dut__.__uuf__._1283_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_112_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2349__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2020_ __dut__._2020_/A1 tie[162] __dut__._2019_/X VGND VGND VPWR VPWR __dut__._3067_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_14_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2922_ clkbuf_5_0_0_tck/X __dut__._2922_/D __dut__._2696_/Y VGND VGND VPWR
+ VPWR __dut__._2922_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2824__CLK __dut__._2846_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1619_ __dut__.__uuf__._1621_/A VGND VGND VPWR VPWR __dut__.__uuf__._1619_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2853_ __dut__._2860_/CLK __dut__._2853_/D __dut__._2765_/Y VGND VGND VPWR
+ VPWR __dut__._2853_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1804_ __dut__._1804_/A1 tie[54] __dut__._1803_/X VGND VGND VPWR VPWR __dut__._2959_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2784_ rst VGND VGND VPWR VPWR __dut__._2784_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1735_ __dut__._2189_/A __dut__._2924_/Q VGND VGND VPWR VPWR __dut__._1735_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_89_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1666_ __dut__._2488_/A1 prod[50] __dut__._1665_/X VGND VGND VPWR VPWR __dut__._2890_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1597_ __dut__._2197_/A __dut__._2854_/Q VGND VGND VPWR VPWR __dut__._1597_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2218_ __dut__._2220_/A1 __dut__._2218_/A2 __dut__._2217_/X VGND VGND VPWR
+ VPWR __dut__._2218_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2149_ __dut__._2207_/A __dut__._2149_/B VGND VGND VPWR VPWR __dut__._2149_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1523__A __dut__.__uuf__._1563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2722__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_169_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2169__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1970_ __dut__.__uuf__._1970_/A VGND VGND VPWR VPWR __dut__.__uuf__._1970_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_23_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1568__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2632__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1404_ __dut__._2315_/B VGND VGND VPWR VPWR __dut__.__uuf__._1404_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_132_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1335_ __dut__.__uuf__._1335_/A VGND VGND VPWR VPWR __dut__.__uuf__._1335_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_120_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1520_ __dut__._1374_/Y mp[10] __dut__._1519_/X VGND VGND VPWR VPWR __dut__._1520_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_116_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1266_ __dut__._2365_/B VGND VGND VPWR VPWR __dut__.__uuf__._1266_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1197_ __dut__.__uuf__._1205_/A VGND VGND VPWR VPWR __dut__.__uuf__._1197_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1451_ __dut__._2509_/A __dut__._2829_/Q VGND VGND VPWR VPWR __dut__._1451_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_74_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1382_ __dut__._1382_/A1 __dut__._1380_/X __dut__._1381_/X VGND VGND VPWR
+ VPWR __dut__._2811_/D sky130_fd_sc_hd__a21o_4
XFILLER_132_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2048__A2 prod[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._3052_ __dut__._3059_/CLK __dut__._3052_/D __dut__._2566_/Y VGND VGND VPWR
+ VPWR __dut__._3052_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2807__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2003_ __dut__._2005_/A __dut__._3058_/Q VGND VGND VPWR VPWR __dut__._2003_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1711__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_261_ _194_/A _261_/D VGND VGND VPWR VPWR _261_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_psn_inst_psn_buff_22_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_192_ _261_/Q _193_/B VGND VGND VPWR VPWR _260_/D sky130_fd_sc_hd__or2_4
XFILLER_50_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2542__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2905_ clkbuf_5_0_0_tck/X __dut__._2905_/D __dut__._2713_/Y VGND VGND VPWR
+ VPWR __dut__._2905_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2836_ __dut__._2836_/CLK __dut__._2836_/D __dut__._2782_/Y VGND VGND VPWR
+ VPWR __dut__._2836_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2767_ rst VGND VGND VPWR VPWR __dut__._2767_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1718_ __dut__._1760_/A1 tie[11] __dut__._1717_/X VGND VGND VPWR VPWR __dut__._2916_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2698_ rst VGND VGND VPWR VPWR __dut__._2698_/Y sky130_fd_sc_hd__inv_2
X__dut__._1649_ __dut__._2491_/A __dut__._2881_/Q VGND VGND VPWR VPWR __dut__._1649_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2717__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_2_0_tck clkbuf_4_3_0_tck/A VGND VGND VPWR VPWR clkbuf_5_5_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_118_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1970__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_286_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1120_ __dut__.__uuf__._1134_/A VGND VGND VPWR VPWR __dut__.__uuf__._1131_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_102_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1051_ __dut__.__uuf__._1214_/A VGND VGND VPWR VPWR __dut__.__uuf__._1051_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2627__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1953_ __dut__.__uuf__._1953_/A VGND VGND VPWR VPWR __dut__.__uuf__._1955_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1531__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1884_ __dut__._1428_/X VGND VGND VPWR VPWR __dut__.__uuf__._1888_/B
+ sky130_fd_sc_hd__inv_2
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2621_ rst VGND VGND VPWR VPWR __dut__._2621_/Y sky130_fd_sc_hd__inv_2
X__dut__._2552_ rst VGND VGND VPWR VPWR __dut__._2552_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2298_ __dut__.__uuf__._2307_/CLK __dut__._2376_/X __dut__.__uuf__._1239_/X
+ VGND VGND VPWR VPWR __dut__._2377_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1318_ __dut__.__uuf__._1335_/A VGND VGND VPWR VPWR __dut__.__uuf__._1318_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_120_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1503_ __dut__._2509_/A __dut__._2842_/Q VGND VGND VPWR VPWR __dut__._1503_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2483_ __dut__._2491_/A prod[50] VGND VGND VPWR VPWR __dut__._2483_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1249_ __dut__.__uuf__._1221_/A __dut__.__uuf__._1248_/Y __dut__.__uuf__._1214_/X
+ __dut__._2373_/B __dut__.__uuf__._1232_/X VGND VGND VPWR VPWR __dut__._2372_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1434_ __dut__._1434_/A1 __dut__._1432_/X __dut__._1433_/X VGND VGND VPWR
+ VPWR __dut__._2824_/D sky130_fd_sc_hd__a21o_4
XFILLER_36_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3104_ __dut__._3106_/CLK __dut__._3104_/D __dut__._2514_/Y VGND VGND VPWR
+ VPWR __dut__._3104_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2537__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3035_ clkbuf_5_4_0_tck/X __dut__._3035_/D __dut__._2583_/Y VGND VGND VPWR
+ VPWR __dut__._3035_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_313_ _313_/CLK _313_/D trst VGND VGND VPWR VPWR _313_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_244_ _312_/Q _311_/Q _244_/C _244_/D VGND VGND VPWR VPWR _244_/X sky130_fd_sc_hd__and4_4
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_175_ _276_/Q _187_/B VGND VGND VPWR VPWR _275_/D sky130_fd_sc_hd__or2_4
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2819_ __dut__._2509_/B __dut__._2819_/D __dut__._2799_/Y VGND VGND VPWR
+ VPWR __dut__._2819_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_111_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3048__CLK __dut__._3058_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2447__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2221_ __dut__.__uuf__._2225_/CLK __dut__._2222_/X __dut__.__uuf__._1576_/X
+ VGND VGND VPWR VPWR __dut__._2223_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_88_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2152_ VGND VGND VPWR VPWR __dut__.__uuf__._2152_/HI tie[159] sky130_fd_sc_hd__conb_1
XFILLER_102_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2083_ VGND VGND VPWR VPWR __dut__.__uuf__._2083_/HI tie[90] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1103_ __dut__.__uuf__._1162_/A VGND VGND VPWR VPWR __dut__.__uuf__._1103_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_84_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1034_ __dut__.__uuf__._1042_/A VGND VGND VPWR VPWR __dut__.__uuf__._1034_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_113_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2357__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1936_ __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR __dut__.__uuf__._1936_/X
+ sky130_fd_sc_hd__buf_2
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1867_ __dut__.__uuf__._1921_/A VGND VGND VPWR VPWR __dut__.__uuf__._1867_/X
+ sky130_fd_sc_hd__buf_2
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1798_ __dut__._2167_/B __dut__._2173_/B VGND VGND VPWR VPWR __dut__.__uuf__._1799_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1983_ __dut__._2005_/A __dut__._3048_/Q VGND VGND VPWR VPWR __dut__._1983_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2604_ rst VGND VGND VPWR VPWR __dut__._2604_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0___dut__.__uuf__.__clk_source__ clkbuf_2_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2535_ rst VGND VGND VPWR VPWR __dut__._2535_/Y sky130_fd_sc_hd__inv_2
X__dut__._2466_ __dut__._2488_/A1 __dut__._2466_/A2 __dut__._2465_/X VGND VGND VPWR
+ VPWR __dut__._2466_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1417_ __dut__._2189_/A __dut__._2819_/Q VGND VGND VPWR VPWR __dut__._1417_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2397_ __dut__._2407_/A prod[7] VGND VGND VPWR VPWR __dut__._2397_/X sky130_fd_sc_hd__and2_4
XFILLER_35_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_5_0___dut__.__uuf__.__clk_source___A clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._3018_ clkbuf_opt_2_tck/A __dut__._3018_/D __dut__._2600_/Y VGND VGND VPWR
+ VPWR __dut__._3018_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_227_ _302_/Q _303_/Q VGND VGND VPWR VPWR _228_/B sky130_fd_sc_hd__or2_4
XFILLER_7_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_158_ _290_/Q _164_/B VGND VGND VPWR VPWR _289_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2730__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2350__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_249_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_151_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2177__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1721_ __dut__.__uuf__._1713_/A __dut__.__uuf__._1718_/B __dut__.__uuf__._1720_/X
+ VGND VGND VPWR VPWR __dut__._2134_/A2 sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1652_ __dut__._1376_/X VGND VGND VPWR VPWR __dut__.__uuf__._1656_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_119_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1583_ __dut__.__uuf__._1584_/A VGND VGND VPWR VPWR __dut__.__uuf__._1583_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_134_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1392__A2 mc[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2640__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2204_ __dut__.__uuf__._2230_/CLK __dut__._2188_/X __dut__.__uuf__._1596_/X
+ VGND VGND VPWR VPWR __dut__._2189_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2135_ VGND VGND VPWR VPWR __dut__.__uuf__._2135_/HI tie[142] sky130_fd_sc_hd__conb_1
XFILLER_130_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2320_ __dut__._2332_/A1 __dut__._2320_/A2 __dut__._2319_/X VGND VGND VPWR
+ VPWR __dut__._2320_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2066_ VGND VGND VPWR VPWR __dut__.__uuf__._2066_/HI tie[73] sky130_fd_sc_hd__conb_1
X__dut__._2251_ __dut__._2251_/A __dut__._2251_/B VGND VGND VPWR VPWR __dut__._2251_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1017_ __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR __dut__.__uuf__._1549_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1616__A __dut__.__uuf__._1628_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2182_ __dut__._2184_/A1 __dut__._2182_/A2 __dut__._2181_/X VGND VGND VPWR
+ VPWR __dut__._2182_/X sky130_fd_sc_hd__a21o_4
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_128 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1876_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_106 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1802_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_117 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1842_/A1 sky130_fd_sc_hd__buf_2
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_139 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2428_/A1 sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1919_ __dut__.__uuf__._1952_/A __dut__.__uuf__._1919_/B __dut__.__uuf__._1919_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1920_/A sky130_fd_sc_hd__or3_4
XFILLER_149_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1966_ __dut__._2004_/A1 tie[135] __dut__._1965_/X VGND VGND VPWR VPWR __dut__._3040_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2550__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1897_ __dut__._2005_/A __dut__._3005_/Q VGND VGND VPWR VPWR __dut__._1897_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2332__A1 __dut__._2332_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2518_ rst VGND VGND VPWR VPWR __dut__._2518_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2449_ __dut__._2507_/A prod[33] VGND VGND VPWR VPWR __dut__._2449_/X sky130_fd_sc_hd__and2_4
XFILLER_35_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2725__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2880__CLK __dut__._3106_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2216__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_131_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__310__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2635__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1704_ __dut__.__uuf__._1982_/A VGND VGND VPWR VPWR __dut__.__uuf__._1704_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1635_ __dut__.__uuf__._1639_/A VGND VGND VPWR VPWR __dut__.__uuf__._1635_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1820_ __dut__._1820_/A1 tie[62] __dut__._1819_/X VGND VGND VPWR VPWR __dut__._2967_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1566_ __dut__.__uuf__._1566_/A VGND VGND VPWR VPWR __dut__.__uuf__._1571_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_150_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1751_ __dut__._2189_/A __dut__._2932_/Q VGND VGND VPWR VPWR __dut__._1751_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1497_ __dut__.__uuf__._1486_/X __dut__.__uuf__._1480_/X __dut__._2273_/B
+ __dut__.__uuf__._1491_/X __dut__.__uuf__._1496_/X VGND VGND VPWR VPWR __dut__._2272_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_135_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1682_ __dut__._2004_/A1 prod[58] __dut__._1681_/X VGND VGND VPWR VPWR __dut__._2898_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2118_ VGND VGND VPWR VPWR __dut__.__uuf__._2118_/HI tie[125] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2049_ VGND VGND VPWR VPWR __dut__.__uuf__._2049_/HI tie[56] sky130_fd_sc_hd__conb_1
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2303_ __dut__._2303_/A __dut__._2303_/B VGND VGND VPWR VPWR __dut__._2303_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3109__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2234_ __dut__._2234_/A1 __dut__._2234_/A2 __dut__._2233_/X VGND VGND VPWR
+ VPWR __dut__._2234_/X sky130_fd_sc_hd__a21o_4
X__dut__._2165_ __dut__._2207_/A __dut__._2165_/B VGND VGND VPWR VPWR __dut__._2165_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2545__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2096_ __dut__._2096_/A1 prod[30] __dut__._2095_/X VGND VGND VPWR VPWR __dut__._3105_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_60_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2239__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_138_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2998_ __dut__._3096_/CLK __dut__._2998_/D __dut__._2620_/Y VGND VGND VPWR
+ VPWR __dut__._2998_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1949_ __dut__._2207_/A __dut__._3031_/Q VGND VGND VPWR VPWR __dut__._1949_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_114_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__145__A3 tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1420_ __dut__.__uuf__._1414_/X __dut__.__uuf__._1419_/X __dut__._2307_/B
+ __dut__.__uuf__._1414_/X VGND VGND VPWR VPWR __dut__._2306_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_156_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1351_ __dut__.__uuf__._1360_/A VGND VGND VPWR VPWR __dut__.__uuf__._1351_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1282_ __dut__.__uuf__._1281_/Y __dut__.__uuf__._1985_/A __dut__.__uuf__._1268_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1282_/X sky130_fd_sc_hd__o21a_4
XFILLER_131_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2365__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2921_ clkbuf_5_0_0_tck/X __dut__._2921_/D __dut__._2697_/Y VGND VGND VPWR
+ VPWR __dut__._2921_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1618_ __dut__.__uuf__._1621_/A VGND VGND VPWR VPWR __dut__.__uuf__._1618_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_107_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2852_ __dut__._2941_/CLK __dut__._2852_/D __dut__._2766_/Y VGND VGND VPWR
+ VPWR __dut__._2852_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1709__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1803_ __dut__._1803_/A __dut__._2958_/Q VGND VGND VPWR VPWR __dut__._1803_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1549_ __dut__.__uuf__._1549_/A VGND VGND VPWR VPWR __dut__.__uuf__._1549_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2783_ rst VGND VGND VPWR VPWR __dut__._2783_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1734_ __dut__._1760_/A1 tie[19] __dut__._1733_/X VGND VGND VPWR VPWR __dut__._2924_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_89_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1665_ __dut__._2491_/A __dut__._2889_/Q VGND VGND VPWR VPWR __dut__._1665_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1596_ __dut__._1374_/Y mc[5] __dut__._1595_/X VGND VGND VPWR VPWR __dut__._1596_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2217_ __dut__._2507_/A __dut__._2217_/B VGND VGND VPWR VPWR __dut__._2217_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_44_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._3081__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2148_ __dut__._2148_/A1 __dut__._2148_/A2 __dut__._2147_/X VGND VGND VPWR
+ VPWR __dut__._2148_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2079_ __dut__._2081_/A __dut__._3096_/Q VGND VGND VPWR VPWR __dut__._2079_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_126_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1619__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_231_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_11_0_tck clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR __dut__._2836_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_36_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2185__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1568__A2 mp[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_26_0_tck clkbuf_5_27_0_tck/A VGND VGND VPWR VPWR _315_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1403_ __dut__.__uuf__._1414_/A VGND VGND VPWR VPWR __dut__.__uuf__._1403_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1334_ __dut__.__uuf__._1327_/X __dut__.__uuf__._1333_/X __dut__._2341_/B
+ __dut__.__uuf__._1327_/X VGND VGND VPWR VPWR __dut__._2340_/A2 sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_4_3_0___dut__.__uuf__.__clk_source__ clkbuf_4_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2293_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1265_ __dut__.__uuf__._1280_/A VGND VGND VPWR VPWR __dut__.__uuf__._1265_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_58_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1196_ __dut__.__uuf__._1192_/X __dut__.__uuf__._1189_/X prod[7]
+ prod[8] __dut__.__uuf__._1185_/X VGND VGND VPWR VPWR __dut__._2396_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1450_ __dut__._1450_/A1 __dut__._1448_/X __dut__._1449_/X VGND VGND VPWR
+ VPWR __dut__._2828_/D sky130_fd_sc_hd__a21o_4
XFILLER_132_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1381_ __dut__._2197_/A __dut__._2874_/Q VGND VGND VPWR VPWR __dut__._1381_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_39_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._3051_ __dut__._3059_/CLK __dut__._3051_/D __dut__._2567_/Y VGND VGND VPWR
+ VPWR __dut__._3051_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2002_ __dut__._2004_/A1 tie[153] __dut__._2001_/X VGND VGND VPWR VPWR __dut__._3058_/D
+ sky130_fd_sc_hd__a21o_4
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_260_ _194_/A _260_/D VGND VGND VPWR VPWR _260_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_191_ _262_/Q _191_/B VGND VGND VPWR VPWR _261_/D sky130_fd_sc_hd__and2_4
XFILLER_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_15_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2904_ __dut__._3079_/CLK __dut__._2904_/D __dut__._2714_/Y VGND VGND VPWR
+ VPWR __dut__._2904_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1439__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2835_ __dut__._2836_/CLK __dut__._2835_/D __dut__._2783_/Y VGND VGND VPWR
+ VPWR __dut__._2835_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2766_ rst VGND VGND VPWR VPWR __dut__._2766_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2697_ rst VGND VGND VPWR VPWR __dut__._2697_/Y sky130_fd_sc_hd__inv_2
X__dut__._1717_ __dut__._2189_/A __dut__._2915_/Q VGND VGND VPWR VPWR __dut__._1717_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_106_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1648_ __dut__._2488_/A1 prod[41] __dut__._1647_/X VGND VGND VPWR VPWR __dut__._2881_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1579_ __dut__._2509_/A __dut__._2861_/Q VGND VGND VPWR VPWR __dut__._1579_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1534__A __dut__.__uuf__._1709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2733__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_279_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1050_ __dut__.__uuf__._1056_/A VGND VGND VPWR VPWR __dut__.__uuf__._1050_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1709__A __dut__.__uuf__._1709_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1952_ __dut__.__uuf__._1952_/A __dut__.__uuf__._1952_/B __dut__.__uuf__._1952_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1953_/A sky130_fd_sc_hd__or3_4
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1883_ __dut__.__uuf__._1875_/A __dut__.__uuf__._1880_/B __dut__.__uuf__._1882_/X
+ VGND VGND VPWR VPWR __dut__._2194_/A2 sky130_fd_sc_hd__o21a_4
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2643__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2620_ rst VGND VGND VPWR VPWR __dut__._2620_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2551_ rst VGND VGND VPWR VPWR __dut__._2551_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2297_ __dut__.__uuf__._2303_/CLK __dut__._2374_/X __dut__.__uuf__._1243_/X
+ VGND VGND VPWR VPWR __dut__._2375_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1317_ __dut__.__uuf__._1311_/X __dut__.__uuf__._1316_/X __dut__._2347_/B
+ __dut__.__uuf__._1311_/X VGND VGND VPWR VPWR __dut__._2346_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1502_ __dut__._1502_/A1 __dut__._1500_/X __dut__._1501_/X VGND VGND VPWR
+ VPWR __dut__._2841_/D sky130_fd_sc_hd__a21o_4
X__dut__._2482_ __dut__._2488_/A1 __dut__._2482_/A2 __dut__._2481_/X VGND VGND VPWR
+ VPWR __dut__._2482_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1248_ __dut__.__uuf__._1248_/A __dut__.__uuf__._1248_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1248_/Y sky130_fd_sc_hd__nand2_4
X__dut__._1433_ __dut__._2507_/A __dut__._2823_/Q VGND VGND VPWR VPWR __dut__._1433_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1179_ __dut__.__uuf__._1208_/A VGND VGND VPWR VPWR __dut__.__uuf__._1191_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_101_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3103_ __dut__._3106_/CLK __dut__._3103_/D __dut__._2515_/Y VGND VGND VPWR
+ VPWR __dut__._3103_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3034_ clkbuf_5_4_0_tck/X __dut__._3034_/D __dut__._2584_/Y VGND VGND VPWR
+ VPWR __dut__._3034_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ _315_/CLK _312_/D trst VGND VGND VPWR VPWR _312_/Q sky130_fd_sc_hd__dfstp_4
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_243_ _301_/Q _300_/Q _302_/Q VGND VGND VPWR VPWR _244_/D sky130_fd_sc_hd__or3_4
XANTENNA___dut__._2553__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_174_ _193_/B VGND VGND VPWR VPWR _187_/B sky130_fd_sc_hd__buf_2
XFILLER_10_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2818_ __dut__._2509_/B __dut__._2818_/D __dut__._2800_/Y VGND VGND VPWR
+ VPWR __dut__._2818_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_3_0_0___dut__.__uuf__.__clk_source___A clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2749_ rst VGND VGND VPWR VPWR __dut__._2749_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2837__CLK __dut__._2846_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1119__A3 prod[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1468__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2728__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2447__B prod[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1640__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2463__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2220_ __dut__.__uuf__._2225_/CLK __dut__._2220_/X __dut__.__uuf__._1577_/X
+ VGND VGND VPWR VPWR __dut__._2221_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_130_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2151_ VGND VGND VPWR VPWR __dut__.__uuf__._2151_/HI tie[158] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2082_ VGND VGND VPWR VPWR __dut__.__uuf__._2082_/HI tie[89] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1102_ __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR __dut__.__uuf__._1162_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_84_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1033_ __dut__.__uuf__._1019_/X __dut__.__uuf__._1023_/X prod[61]
+ prod[62] __dut__.__uuf__._1025_/X VGND VGND VPWR VPWR __dut__._2504_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_110_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2638__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1935_ __dut__.__uuf__._1935_/A VGND VGND VPWR VPWR __dut__._2216_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1866_ __dut__.__uuf__._1866_/A VGND VGND VPWR VPWR __dut__.__uuf__._1869_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_138_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1797_ __dut__._1392_/X VGND VGND VPWR VPWR __dut__.__uuf__._1801_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2373__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1982_ __dut__._2004_/A1 tie[143] __dut__._1981_/X VGND VGND VPWR VPWR __dut__._3048_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_138_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2272__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_152_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2603_ rst VGND VGND VPWR VPWR __dut__._2603_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2349_ __dut__.__uuf__._2353_/CLK __dut__._2478_/X __dut__.__uuf__._1071_/X
+ VGND VGND VPWR VPWR prod[48] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1717__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_1_0_tck clkbuf_4_1_0_tck/A VGND VGND VPWR VPWR clkbuf_5_3_0_tck/A sky130_fd_sc_hd__clkbuf_1
X__dut__._2534_ rst VGND VGND VPWR VPWR __dut__._2534_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_82_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2465_ __dut__._2491_/A prod[41] VGND VGND VPWR VPWR __dut__._2465_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2548__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1416_ __dut__._1374_/Y mc[19] __dut__._1415_/X VGND VGND VPWR VPWR __dut__._1416_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._2396_ __dut__._2412_/A1 __dut__._2396_/A2 __dut__._2395_/X VGND VGND VPWR
+ VPWR __dut__._2396_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3017_ clkbuf_5_6_0_tck/X __dut__._3017_/D __dut__._2601_/Y VGND VGND VPWR
+ VPWR __dut__._3017_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1037__A2 __dut__.__uuf__._1023_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_226_ _301_/Q _300_/Q _222_/A VGND VGND VPWR VPWR _300_/D sky130_fd_sc_hd__o21a_4
X_157_ tdi _164_/B VGND VGND VPWR VPWR _290_/D sky130_fd_sc_hd__and2_4
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1627__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3015__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2102__A2 prod[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_144_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1720_ __dut__.__uuf__._1828_/A VGND VGND VPWR VPWR __dut__.__uuf__._1720_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1651_ __dut__.__uuf__._1904_/A VGND VGND VPWR VPWR __dut__.__uuf__._1680_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1582_ __dut__.__uuf__._1584_/A VGND VGND VPWR VPWR __dut__.__uuf__._1582_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_134_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2203_ __dut__.__uuf__._2240_/CLK __dut__._2186_/X __dut__.__uuf__._1598_/X
+ VGND VGND VPWR VPWR __dut__._2187_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2134_ VGND VGND VPWR VPWR __dut__.__uuf__._2134_/HI tie[141] sky130_fd_sc_hd__conb_1
XFILLER_130_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2065_ VGND VGND VPWR VPWR __dut__.__uuf__._2065_/HI tie[72] sky130_fd_sc_hd__conb_1
XFILLER_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2250_ __dut__._2250_/A1 __dut__._2250_/A2 __dut__._2249_/X VGND VGND VPWR
+ VPWR __dut__._2250_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1016_ __dut__.__uuf__._1989_/A __dut__._2109_/B __dut__.__uuf__._1016_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1176_/A sky130_fd_sc_hd__or3_4
XFILLER_72_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2181_ __dut__._2189_/A __dut__._2181_/B VGND VGND VPWR VPWR __dut__._2181_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_140_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_107 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1804_/A1 sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1604__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_118 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1844_/A1 sky130_fd_sc_hd__buf_2
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_129 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1878_/A1 sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1918_ __dut__._2211_/B __dut__._2217_/B __dut__.__uuf__._1917_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1919_/C sky130_fd_sc_hd__o21ai_4
XFILLER_149_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1849_ __dut__.__uuf__._1842_/A __dut__.__uuf__._1847_/B __dut__.__uuf__._1828_/X
+ VGND VGND VPWR VPWR __dut__._2182_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1965_ __dut__._1965_/A __dut__._3039_/Q VGND VGND VPWR VPWR __dut__._1965_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_4_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1896_ __dut__._2004_/A1 tie[100] __dut__._1895_/X VGND VGND VPWR VPWR __dut__._3005_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1447__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2517_ rst VGND VGND VPWR VPWR __dut__._2517_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2168__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2448_ __dut__._2448_/A1 __dut__._2448_/A2 __dut__._2447_/X VGND VGND VPWR
+ VPWR __dut__._2448_/X sky130_fd_sc_hd__a21o_4
XFILLER_114_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2379_ __dut__._2407_/A __dut__._2379_/B VGND VGND VPWR VPWR __dut__._2379_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_90_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_209_ _247_/Q VGND VGND VPWR VPWR _209_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2741__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_261_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1703_ __dut__.__uuf__._1703_/A VGND VGND VPWR VPWR __dut__.__uuf__._1982_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1634_ __dut__.__uuf__._1640_/A VGND VGND VPWR VPWR __dut__.__uuf__._1639_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2651__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1565_ __dut__.__uuf__._1549_/X __dut__.__uuf__._1828_/A __dut__._2239_/B
+ __dut__.__uuf__._1447_/A __dut__.__uuf__._1564_/X VGND VGND VPWR VPWR __dut__._2238_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_135_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1750_ __dut__._1760_/A1 tie[27] __dut__._1749_/X VGND VGND VPWR VPWR __dut__._2932_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_150_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1496_ __dut__._1548_/X __dut__.__uuf__._1487_/X __dut__._2275_/B
+ __dut__.__uuf__._1492_/X VGND VGND VPWR VPWR __dut__.__uuf__._1496_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1681_ __dut__._1891_/A __dut__._2897_/Q VGND VGND VPWR VPWR __dut__._1681_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_142_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2117_ VGND VGND VPWR VPWR __dut__.__uuf__._2117_/HI tie[124] sky130_fd_sc_hd__conb_1
XFILLER_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._2048_ VGND VGND VPWR VPWR __dut__.__uuf__._2048_/HI tie[55] sky130_fd_sc_hd__conb_1
X__dut__._2302_ __dut__._2308_/A1 __dut__._2302_/A2 __dut__._2301_/X VGND VGND VPWR
+ VPWR __dut__._2302_/X sky130_fd_sc_hd__a21o_4
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2233_ __dut__._2325_/A __dut__._2233_/B VGND VGND VPWR VPWR __dut__._2233_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2164_ __dut__._2172_/A1 __dut__._2164_/A2 __dut__._2163_/X VGND VGND VPWR
+ VPWR __dut__._2164_/X sky130_fd_sc_hd__a21o_4
XFILLER_25_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_45_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2095_ __dut__._2095_/A __dut__._3104_/Q VGND VGND VPWR VPWR __dut__._2095_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2002__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2561__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2997_ __dut__._3096_/CLK __dut__._2997_/D __dut__._2621_/Y VGND VGND VPWR
+ VPWR __dut__._2997_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1948_ __dut__._2172_/A1 tie[126] __dut__._1947_/X VGND VGND VPWR VPWR __dut__._3031_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1879_ __dut__._1881_/A __dut__._2996_/Q VGND VGND VPWR VPWR __dut__._1879_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1905__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__271__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2736__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2455__B prod[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_107_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2471__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1350_ __dut__.__uuf__._1338_/X __dut__.__uuf__._1349_/X __dut__._2335_/B
+ __dut__.__uuf__._1338_/X VGND VGND VPWR VPWR __dut__._2334_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1281_ __dut__._2361_/B VGND VGND VPWR VPWR __dut__.__uuf__._1281_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_124_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2480__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2646__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2920_ clkbuf_5_0_0_tck/X __dut__._2920_/D __dut__._2698_/Y VGND VGND VPWR
+ VPWR __dut__._2920_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2851_ __dut__._2941_/CLK __dut__._2851_/D __dut__._2767_/Y VGND VGND VPWR
+ VPWR __dut__._2851_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2381__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1617_ __dut__.__uuf__._1621_/A VGND VGND VPWR VPWR __dut__.__uuf__._1617_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1802_ __dut__._1802_/A1 tie[53] __dut__._1801_/X VGND VGND VPWR VPWR __dut__._2958_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_146_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1548_ __dut__.__uuf__._1562_/A VGND VGND VPWR VPWR __dut__.__uuf__._1548_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2782_ rst VGND VGND VPWR VPWR __dut__._2782_/Y sky130_fd_sc_hd__inv_2
X__dut__._1733_ __dut__._2189_/A __dut__._2923_/Q VGND VGND VPWR VPWR __dut__._1733_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1479_ __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR __dut__.__uuf__._1479_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_103_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1664_ __dut__._2488_/A1 prod[49] __dut__._1663_/X VGND VGND VPWR VPWR __dut__._2889_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_131_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1725__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1595_ __dut__._2509_/A __dut__._2865_/Q VGND VGND VPWR VPWR __dut__._1595_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_85_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2206__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2216_ __dut__._2220_/A1 __dut__._2216_/A2 __dut__._2215_/X VGND VGND VPWR
+ VPWR __dut__._2216_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2556__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2147_ __dut__._2207_/A __dut__._2147_/B VGND VGND VPWR VPWR __dut__._2147_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2078_ __dut__._2078_/A1 prod[21] __dut__._2077_/X VGND VGND VPWR VPWR __dut__._3096_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_145_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_224_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2462__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_290 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1797_/A sky130_fd_sc_hd__buf_2
XFILLER_145_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1402_ __dut__.__uuf__._1411_/A VGND VGND VPWR VPWR __dut__.__uuf__._1402_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_144_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1333_ __dut__.__uuf__._1332_/Y __dut__.__uuf__._1321_/X __dut__.__uuf__._1322_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1333_/X sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._2893__CLK __dut__._3106_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1264_ __dut__.__uuf__._1261_/X __dut__.__uuf__._1988_/B __dut__._2239_/B
+ __dut__.__uuf__._1025_/X VGND VGND VPWR VPWR __dut__._2366_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1195_ __dut__.__uuf__._1205_/A VGND VGND VPWR VPWR __dut__.__uuf__._1195_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1177__A __dut__.__uuf__._1463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1560__B2 __dut__.__uuf__._1294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1380_ __dut__._1374_/Y mc[10] __dut__._1379_/X VGND VGND VPWR VPWR __dut__._1380_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2229__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_67_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3050_ __dut__._3058_/CLK __dut__._3050_/D __dut__._2568_/Y VGND VGND VPWR
+ VPWR __dut__._3050_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2001_ __dut__._2005_/A __dut__._3057_/Q VGND VGND VPWR VPWR __dut__._2001_/X
+ sky130_fd_sc_hd__and2_4
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_190_ _263_/Q _191_/B VGND VGND VPWR VPWR _262_/D sky130_fd_sc_hd__and2_4
XFILLER_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1640__A __dut__.__uuf__._1640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2903_ __dut__._3079_/CLK __dut__._2903_/D __dut__._2715_/Y VGND VGND VPWR
+ VPWR __dut__._2903_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2834_ __dut__._2836_/CLK __dut__._2834_/D __dut__._2784_/Y VGND VGND VPWR
+ VPWR __dut__._2834_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2765_ rst VGND VGND VPWR VPWR __dut__._2765_/Y sky130_fd_sc_hd__inv_2
X__dut__._1716_ __dut__._1760_/A1 tie[10] __dut__._1715_/X VGND VGND VPWR VPWR __dut__._2915_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_150_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2696_ rst VGND VGND VPWR VPWR __dut__._2696_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1455__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1647_ __dut__._2491_/A __dut__._2880_/Q VGND VGND VPWR VPWR __dut__._1647_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1578_ __dut__._1780_/A1 __dut__._1576_/X __dut__._1577_/X VGND VGND VPWR
+ VPWR __dut__._2860_/D sky130_fd_sc_hd__a21o_4
XFILLER_64_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_13_0___dut__.__uuf__.__clk_source__ clkbuf_3_6_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2288_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_122_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0___dut__.__uuf__.__clk_source__ __dut__._2510_/X VGND VGND VPWR VPWR clkbuf_0___dut__.__uuf__.__clk_source__/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_174_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1951_ __dut__._2223_/B __dut__._2229_/B __dut__.__uuf__._1950_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1952_/C sky130_fd_sc_hd__o21ai_4
X__dut__.__uuf__._1882_ __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR __dut__.__uuf__._1882_/X
+ sky130_fd_sc_hd__buf_2
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1316_ __dut__.__uuf__._1315_/Y __dut__.__uuf__._1294_/X __dut__.__uuf__._1296_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1316_/X sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._3071__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2550_ rst VGND VGND VPWR VPWR __dut__._2550_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2296_ __dut__.__uuf__._2303_/CLK __dut__._2372_/X __dut__.__uuf__._1247_/X
+ VGND VGND VPWR VPWR __dut__._2373_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_143_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1501_ __dut__._2189_/A __dut__._2840_/Q VGND VGND VPWR VPWR __dut__._1501_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2481_ __dut__._2491_/A prod[49] VGND VGND VPWR VPWR __dut__._2481_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1247_ __dut__.__uuf__._1254_/A VGND VGND VPWR VPWR __dut__.__uuf__._1247_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1432_ __dut__._1374_/Y mc[22] __dut__._1431_/X VGND VGND VPWR VPWR __dut__._1432_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1178_ __dut__.__uuf__._1177_/X __dut__.__uuf__._1173_/X prod[13]
+ prod[14] __dut__.__uuf__._1170_/X VGND VGND VPWR VPWR __dut__._2408_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._3102_ __dut__._3102_/CLK __dut__._3102_/D __dut__._2516_/Y VGND VGND VPWR
+ VPWR __dut__._3102_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3033_ clkbuf_5_1_0_tck/X __dut__._3033_/D __dut__._2585_/Y VGND VGND VPWR
+ VPWR __dut__._3033_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_311_ _315_/CLK _311_/D trst VGND VGND VPWR VPWR _311_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1049__B1 prod[57] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_242_ _242_/A VGND VGND VPWR VPWR _244_/C sky130_fd_sc_hd__inv_2
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_173_ _277_/Q _173_/B VGND VGND VPWR VPWR _276_/D sky130_fd_sc_hd__and2_4
XFILLER_10_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2817_ __dut__._2509_/B __dut__._2817_/D __dut__._2801_/Y VGND VGND VPWR
+ VPWR __dut__._2817_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_5_10_0_tck clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR __dut__._2846_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_151_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2748_ rst VGND VGND VPWR VPWR __dut__._2748_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2679_ rst VGND VGND VPWR VPWR __dut__._2679_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_25_0_tck clkbuf_5_25_0_tck/A VGND VGND VPWR VPWR _290_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1468__A2 mc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1913__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1640__A2 prod[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2744__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_291_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__304__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2150_ VGND VGND VPWR VPWR __dut__.__uuf__._2150_/HI tie[157] sky130_fd_sc_hd__conb_1
XFILLER_88_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2081_ VGND VGND VPWR VPWR __dut__.__uuf__._2081_/HI tie[88] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1101_ __dut__.__uuf__._1101_/A VGND VGND VPWR VPWR __dut__.__uuf__._1101_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1032_ __dut__.__uuf__._1042_/A VGND VGND VPWR VPWR __dut__.__uuf__._1032_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_110_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1823__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2408__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1934_ __dut__.__uuf__._1975_/A __dut__.__uuf__._1934_/B __dut__.__uuf__._1934_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1935_/A sky130_fd_sc_hd__or3_4
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2654__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1865_ __dut__.__uuf__._1898_/A __dut__.__uuf__._1865_/B __dut__.__uuf__._1865_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1866_/A sky130_fd_sc_hd__or3_4
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1796_ __dut__.__uuf__._1904_/A VGND VGND VPWR VPWR __dut__.__uuf__._1844_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_149_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1981_ __dut__._2005_/A __dut__._3047_/Q VGND VGND VPWR VPWR __dut__._1981_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_138_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2602_ rst VGND VGND VPWR VPWR __dut__._2602_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2348_ __dut__.__uuf__._2353_/CLK __dut__._2476_/X __dut__.__uuf__._1077_/X
+ VGND VGND VPWR VPWR prod[47] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2279_ __dut__.__uuf__._2288_/CLK __dut__._2338_/X __dut__.__uuf__._1335_/X
+ VGND VGND VPWR VPWR __dut__._2339_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2533_ rst VGND VGND VPWR VPWR __dut__._2533_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1733__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2464_ __dut__._2488_/A1 __dut__._2464_/A2 __dut__._2463_/X VGND VGND VPWR
+ VPWR __dut__._2464_/X sky130_fd_sc_hd__a21o_4
XFILLER_62_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_75_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1415_ __dut__._2509_/A __dut__._2820_/Q VGND VGND VPWR VPWR __dut__._1415_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2395_ __dut__._2407_/A prod[6] VGND VGND VPWR VPWR __dut__._2395_/X sky130_fd_sc_hd__and2_4
XFILLER_103_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3016_ clkbuf_5_5_0_tck/X __dut__._3016_/D __dut__._2602_/Y VGND VGND VPWR
+ VPWR __dut__._3016_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2564__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1037__A3 prod[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_225_ _300_/Q _225_/B VGND VGND VPWR VPWR _299_/D sky130_fd_sc_hd__and2_4
XFILLER_143_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_156_ _183_/A VGND VGND VPWR VPWR _164_/B sky130_fd_sc_hd__buf_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2739__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_137_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1650_ __dut__.__uuf__._1703_/A VGND VGND VPWR VPWR __dut__.__uuf__._1904_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_147_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1581_ __dut__.__uuf__._1584_/A VGND VGND VPWR VPWR __dut__.__uuf__._1581_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_146_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2202_ __dut__.__uuf__._2240_/CLK __dut__._2184_/X __dut__.__uuf__._1599_/X
+ VGND VGND VPWR VPWR __dut__._2185_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2133_ VGND VGND VPWR VPWR __dut__.__uuf__._2133_/HI tie[140] sky130_fd_sc_hd__conb_1
XFILLER_88_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2649__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2064_ VGND VGND VPWR VPWR __dut__.__uuf__._2064_/HI tie[71] sky130_fd_sc_hd__conb_1
XFILLER_84_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1015_ __dut__.__uuf__._1989_/C VGND VGND VPWR VPWR __dut__.__uuf__._1016_/C
+ sky130_fd_sc_hd__inv_2
XFILLER_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2180_ __dut__._2184_/A1 __dut__._2180_/A2 __dut__._2179_/X VGND VGND VPWR
+ VPWR __dut__._2180_/X sky130_fd_sc_hd__a21o_4
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_108 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1806_/A1 sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1604__A2 mp[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_119 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._2044_/A1 sky130_fd_sc_hd__buf_2
XFILLER_25_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__297__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1917_ __dut__.__uuf__._1917_/A VGND VGND VPWR VPWR __dut__.__uuf__._1917_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1848_ __dut__.__uuf__._1848_/A VGND VGND VPWR VPWR __dut__._2184_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_138_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1779_ __dut__._2159_/B __dut__._2165_/B __dut__.__uuf__._1778_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1780_/C sky130_fd_sc_hd__o21ai_4
XFILLER_126_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1964_ __dut__._2004_/A1 tie[134] __dut__._1963_/X VGND VGND VPWR VPWR __dut__._3039_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_153_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1895_ __dut__._2005_/A __dut__._3004_/Q VGND VGND VPWR VPWR __dut__._1895_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1540__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2559__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2516_ rst VGND VGND VPWR VPWR __dut__._2516_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_9_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2447_ __dut__._2507_/A prod[32] VGND VGND VPWR VPWR __dut__._2447_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1463__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2378_ __dut__._2412_/A1 __dut__._2378_/A2 __dut__._2377_/X VGND VGND VPWR
+ VPWR __dut__._2378_/X sky130_fd_sc_hd__a21o_4
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_208_ _252_/Q _208_/B VGND VGND VPWR VPWR _208_/X sky130_fd_sc_hd__or2_4
XFILLER_156_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_139_ _238_/B _138_/B _138_/Y _128_/X VGND VGND VPWR VPWR _140_/A sky130_fd_sc_hd__a211o_4
XFILLER_124_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2469__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_254_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1373__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1702_ __dut__.__uuf__._1702_/A VGND VGND VPWR VPWR __dut__.__uuf__._1706_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1633_ __dut__.__uuf__._1633_/A VGND VGND VPWR VPWR __dut__.__uuf__._1633_/X
+ sky130_fd_sc_hd__buf_2
Xclkbuf_4_0_0_tck clkbuf_4_1_0_tck/A VGND VGND VPWR VPWR clkbuf_5_1_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1564_ __dut__._1476_/X __dut__.__uuf__._1550_/X __dut__._2241_/B
+ __dut__.__uuf__._1294_/A VGND VGND VPWR VPWR __dut__.__uuf__._1564_/X sky130_fd_sc_hd__o22a_4
XFILLER_135_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1495_ __dut__.__uuf__._1501_/A VGND VGND VPWR VPWR __dut__.__uuf__._1495_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1680_ __dut__._2502_/A1 prod[57] __dut__._1679_/X VGND VGND VPWR VPWR __dut__._2897_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2116_ VGND VGND VPWR VPWR __dut__.__uuf__._2116_/HI tie[123] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2379__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2047_ VGND VGND VPWR VPWR __dut__.__uuf__._2047_/HI tie[54] sky130_fd_sc_hd__conb_1
X__dut__._2301_ __dut__._2303_/A __dut__._2301_/B VGND VGND VPWR VPWR __dut__._2301_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2232_ __dut__._2232_/A1 __dut__._2232_/A2 __dut__._2231_/X VGND VGND VPWR
+ VPWR __dut__._2232_/X sky130_fd_sc_hd__a21o_4
XFILLER_84_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2163_ __dut__._2207_/A __dut__._2163_/B VGND VGND VPWR VPWR __dut__._2163_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2094_ __dut__._2094_/A1 prod[29] __dut__._2093_/X VGND VGND VPWR VPWR __dut__._3104_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_80_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_38_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2996_ __dut__._3096_/CLK __dut__._2996_/D __dut__._2622_/Y VGND VGND VPWR
+ VPWR __dut__._2996_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1947_ __dut__._2207_/A __dut__._3030_/Q VGND VGND VPWR VPWR __dut__._1947_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_140_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1878_ __dut__._1878_/A1 tie[91] __dut__._1877_/X VGND VGND VPWR VPWR __dut__._2996_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_121_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1921__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2752__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1504__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1280_ __dut__.__uuf__._1280_/A VGND VGND VPWR VPWR __dut__.__uuf__._1280_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2199__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1831__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3028__CLK clkbuf_5_1_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1463__A __dut__.__uuf__._1463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2662__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1616_ __dut__.__uuf__._1628_/A VGND VGND VPWR VPWR __dut__.__uuf__._1621_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._2850_ __dut__._2941_/CLK __dut__._2850_/D __dut__._2768_/Y VGND VGND VPWR
+ VPWR __dut__._2850_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1801_ __dut__._1801_/A __dut__._2957_/Q VGND VGND VPWR VPWR __dut__._1801_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1547_ __dut__.__uuf__._1566_/A VGND VGND VPWR VPWR __dut__.__uuf__._1562_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._2781_ rst VGND VGND VPWR VPWR __dut__._2781_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1732_ __dut__._1760_/A1 tie[18] __dut__._1731_/X VGND VGND VPWR VPWR __dut__._2923_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1478_ __dut__.__uuf__._1463_/X __dut__.__uuf__._1458_/X __dut__._2281_/B
+ __dut__.__uuf__._1469_/X __dut__.__uuf__._1477_/X VGND VGND VPWR VPWR __dut__._2280_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_150_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1663_ __dut__._2491_/A __dut__._2888_/Q VGND VGND VPWR VPWR __dut__._1663_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_131_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1594_ __dut__._1780_/A1 __dut__._1592_/X __dut__._1593_/X VGND VGND VPWR
+ VPWR __dut__._2864_/D sky130_fd_sc_hd__a21o_4
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1741__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2215_ __dut__._2507_/A __dut__._2215_/B VGND VGND VPWR VPWR __dut__._2215_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2146_ __dut__._2148_/A1 __dut__._2146_/A2 __dut__._2145_/X VGND VGND VPWR
+ VPWR __dut__._2146_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_7_0_tck clkbuf_3_7_0_tck/A VGND VGND VPWR VPWR clkbuf_3_7_0_tck/X sky130_fd_sc_hd__clkbuf_1
X__dut__._2077_ __dut__._2081_/A __dut__._3095_/Q VGND VGND VPWR VPWR __dut__._2077_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1982__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2572__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2979_ __dut__._3079_/CLK __dut__._2979_/D __dut__._2639_/Y VGND VGND VPWR
+ VPWR __dut__._2979_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_141_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2747__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1651__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_217_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2300__CLK __dut__.__uuf__._2303_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_31_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpsn_inst_psn_buff_280 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2325_/A sky130_fd_sc_hd__buf_4
Xpsn_inst_psn_buff_291 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1821_/A sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1401_ __dut__.__uuf__._1389_/X __dut__.__uuf__._1400_/X __dut__._2315_/B
+ __dut__.__uuf__._1389_/X VGND VGND VPWR VPWR __dut__._2314_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1332_ __dut__._2343_/B VGND VGND VPWR VPWR __dut__.__uuf__._1332_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_132_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1263_ __dut__.__uuf__._1533_/A VGND VGND VPWR VPWR __dut__.__uuf__._1988_/B
+ sky130_fd_sc_hd__buf_2
XFILLER_113_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1458__A __dut__.__uuf__._1480_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1194_ __dut__.__uuf__._1208_/A VGND VGND VPWR VPWR __dut__.__uuf__._1205_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_86_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2657__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2000_ __dut__._2004_/A1 tie[152] __dut__._1999_/X VGND VGND VPWR VPWR __dut__._3057_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_42_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1964__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2902_ __dut__._3109_/CLK __dut__._2902_/D __dut__._2716_/Y VGND VGND VPWR
+ VPWR __dut__._2902_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2833_ __dut__._2860_/CLK __dut__._2833_/D __dut__._2785_/Y VGND VGND VPWR
+ VPWR __dut__._2833_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2764_ rst VGND VGND VPWR VPWR __dut__._2764_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1715_ __dut__._2189_/A __dut__._2914_/Q VGND VGND VPWR VPWR __dut__._1715_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2695_ rst VGND VGND VPWR VPWR __dut__._2695_/Y sky130_fd_sc_hd__inv_2
X__dut__._1646_ __dut__._2502_/A1 prod[40] __dut__._1645_/X VGND VGND VPWR VPWR __dut__._2880_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1577_ __dut__._1589_/A __dut__._2859_/Q VGND VGND VPWR VPWR __dut__._1577_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2567__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1471__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0___dut__.__uuf__.__clk_source__/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2129_ __dut__._2141_/A __dut__._2129_/B VGND VGND VPWR VPWR __dut__._2129_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_146_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2380__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_167_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2477__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1950_ __dut__.__uuf__._1950_/A VGND VGND VPWR VPWR __dut__.__uuf__._1950_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1881_ __dut__.__uuf__._1881_/A VGND VGND VPWR VPWR __dut__._2196_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_23_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__284__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1946__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2860__CLK __dut__._2860_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2364_ __dut__.__uuf__._2364_/CLK __dut__._2508_/X __dut__.__uuf__._1992_/X
+ VGND VGND VPWR VPWR prod[63] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1315_ __dut__._2349_/B VGND VGND VPWR VPWR __dut__.__uuf__._1315_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1188__A __dut__.__uuf__._1464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2295_ __dut__.__uuf__._2307_/CLK __dut__._2370_/X __dut__.__uuf__._1250_/X
+ VGND VGND VPWR VPWR __dut__._2371_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_143_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2480_ __dut__._2488_/A1 __dut__._2480_/A2 __dut__._2479_/X VGND VGND VPWR
+ VPWR __dut__._2480_/X sky130_fd_sc_hd__a21o_4
X__dut__._1500_ __dut__._1374_/Y mp[6] __dut__._1499_/X VGND VGND VPWR VPWR __dut__._1500_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1246_ __dut__.__uuf__._1244_/Y __dut__.__uuf__._1245_/X __dut__.__uuf__._1214_/X
+ __dut__._2375_/B __dut__.__uuf__._1232_/X VGND VGND VPWR VPWR __dut__._2374_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_47_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1431_ __dut__._2509_/A __dut__._2824_/Q VGND VGND VPWR VPWR __dut__._1431_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1177_ __dut__.__uuf__._1463_/A VGND VGND VPWR VPWR __dut__.__uuf__._1177_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3101_ __dut__._3102_/CLK __dut__._3101_/D __dut__._2517_/Y VGND VGND VPWR
+ VPWR __dut__._3101_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_310_ _315_/CLK _310_/D trst VGND VGND VPWR VPWR _310_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._3032_ clkbuf_5_1_0_tck/X __dut__._3032_/D __dut__._2586_/Y VGND VGND VPWR
+ VPWR __dut__._3032_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1651__A __dut__.__uuf__._1904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_241_ tms _240_/X _128_/X VGND VGND VPWR VPWR _306_/D sky130_fd_sc_hd__a21o_4
XFILLER_156_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_psn_inst_psn_buff_20_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_172_ _278_/Q _172_/B VGND VGND VPWR VPWR _277_/D sky130_fd_sc_hd__or2_4
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._2816_ __dut__._2509_/B __dut__._2816_/D __dut__._2802_/Y VGND VGND VPWR
+ VPWR __dut__._2816_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2362__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2747_ rst VGND VGND VPWR VPWR __dut__._2747_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2678_ rst VGND VGND VPWR VPWR __dut__._2678_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1629_ __dut__._2197_/A __dut__._2872_/Q VGND VGND VPWR VPWR __dut__._1629_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2883__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2760__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1212__A1 __dut__.__uuf__._1206_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_284_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1100_ __dut__.__uuf__._1088_/X __dut__.__uuf__._1099_/X prod[39]
+ prod[40] __dut__.__uuf__._1096_/X VGND VGND VPWR VPWR __dut__._2460_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._2080_ VGND VGND VPWR VPWR __dut__.__uuf__._2080_/HI tie[87] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1031_ __dut__.__uuf__._1019_/X __dut__.__uuf__._1023_/X prod[62]
+ prod[63] __dut__.__uuf__._1025_/X VGND VGND VPWR VPWR __dut__._2506_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1933_ __dut__.__uuf__._1921_/X __dut__.__uuf__._1931_/B __dut__.__uuf__._1931_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1934_/C sky130_fd_sc_hd__o21a_4
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1864_ __dut__._2191_/B __dut__._2197_/B __dut__.__uuf__._1863_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1865_/C sky130_fd_sc_hd__o21ai_4
X__dut__.__uuf__._1795_ __dut__.__uuf__._1788_/A __dut__.__uuf__._1793_/B __dut__.__uuf__._1774_/X
+ VGND VGND VPWR VPWR __dut__._2162_/A2 sky130_fd_sc_hd__o21a_4
X__dut__._1980_ __dut__._2004_/A1 tie[142] __dut__._1979_/X VGND VGND VPWR VPWR __dut__._3047_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_138_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2670__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2344__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2601_ rst VGND VGND VPWR VPWR __dut__._2601_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2347_ __dut__.__uuf__._2353_/CLK __dut__._2474_/X __dut__.__uuf__._1079_/X
+ VGND VGND VPWR VPWR prod[46] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2532_ rst VGND VGND VPWR VPWR __dut__._2532_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2278_ __dut__.__uuf__._2278_/CLK __dut__._2336_/X __dut__.__uuf__._1341_/X
+ VGND VGND VPWR VPWR __dut__._2337_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1229_ __dut__.__uuf__._1229_/A __dut__.__uuf__._1292_/A VGND VGND
+ VPWR VPWR __dut__.__uuf__._1446_/A sky130_fd_sc_hd__or2_4
XFILLER_87_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2463_ __dut__._2491_/A prod[40] VGND VGND VPWR VPWR __dut__._2463_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1646__A __dut__.__uuf__._1992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1414_ __dut__._1414_/A1 __dut__._1412_/X __dut__._1413_/X VGND VGND VPWR
+ VPWR __dut__._2819_/D sky130_fd_sc_hd__a21o_4
X__dut__._2394_ __dut__._2412_/A1 __dut__._2394_/A2 __dut__._2393_/X VGND VGND VPWR
+ VPWR __dut__._2394_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_68_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._3015_ clkbuf_5_5_0_tck/X __dut__._3015_/D __dut__._2603_/Y VGND VGND VPWR
+ VPWR __dut__._3015_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_224_ _301_/Q _299_/Q _232_/A VGND VGND VPWR VPWR _298_/D sky130_fd_sc_hd__o21a_4
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_155_ _193_/B VGND VGND VPWR VPWR _183_/A sky130_fd_sc_hd__inv_2
XFILLER_6_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2580__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2755__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3061__CLK clkbuf_5_6_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1580_ __dut__.__uuf__._1584_/A VGND VGND VPWR VPWR __dut__.__uuf__._1580_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_146_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2326__A1 __dut__._2332_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2191__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_108_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2201_ __dut__.__uuf__._2240_/CLK __dut__._2182_/X __dut__.__uuf__._1600_/X
+ VGND VGND VPWR VPWR __dut__._2183_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_142_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2132_ VGND VGND VPWR VPWR __dut__.__uuf__._2132_/HI tie[139] sky130_fd_sc_hd__conb_1
XFILLER_115_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2063_ VGND VGND VPWR VPWR __dut__.__uuf__._2063_/HI tie[70] sky130_fd_sc_hd__conb_1
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1014_ __dut__._2373_/B __dut__.__uuf__._1219_/A __dut__._2369_/B
+ __dut__.__uuf__._1014_/D VGND VGND VPWR VPWR __dut__.__uuf__._1989_/C sky130_fd_sc_hd__or4_4
XFILLER_29_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__.__uuf__._1672__A1 __dut__.__uuf__._1261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_109 __dut__._1418_/A1 VGND VGND VPWR VPWR __dut__._1818_/A1 sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2665__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1916_ __dut__._2211_/B __dut__._2217_/B VGND VGND VPWR VPWR __dut__.__uuf__._1917_/A
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1847_ __dut__.__uuf__._1869_/A __dut__.__uuf__._1847_/B __dut__.__uuf__._1847_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1848_/A sky130_fd_sc_hd__or3_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_24_0_tck clkbuf_5_25_0_tck/A VGND VGND VPWR VPWR _313_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_20_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1778_ __dut__.__uuf__._1778_/A VGND VGND VPWR VPWR __dut__.__uuf__._1778_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_125_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1963_ __dut__._1963_/A __dut__._3038_/Q VGND VGND VPWR VPWR __dut__._1963_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_146_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1894_ __dut__._2004_/A1 tie[99] __dut__._1893_/X VGND VGND VPWR VPWR __dut__._3004_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_121_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1540__A2 mp[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2515_ rst VGND VGND VPWR VPWR __dut__._2515_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2446_ __dut__._2446_/A1 __dut__._2446_/A2 __dut__._2445_/X VGND VGND VPWR
+ VPWR __dut__._2446_/X sky130_fd_sc_hd__a21o_4
XFILLER_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1112__B1 prod[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2377_ __dut__._2407_/A __dut__._2377_/B VGND VGND VPWR VPWR __dut__._2377_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._3084__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2575__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1919__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_207_ _211_/A VGND VGND VPWR VPWR _208_/B sky130_fd_sc_hd__inv_2
XFILLER_144_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_138_ _307_/Q _138_/B VGND VGND VPWR VPWR _138_/Y sky130_fd_sc_hd__nor2_4
XFILLER_143_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_247_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2485__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1701_ __dut__.__uuf__._1736_/A __dut__.__uuf__._1701_/B __dut__.__uuf__._1701_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1702_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1632_ __dut__.__uuf__._1633_/A VGND VGND VPWR VPWR __dut__.__uuf__._1632_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_119_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1563_ __dut__.__uuf__._1563_/A VGND VGND VPWR VPWR __dut__.__uuf__._1828_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_128_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1494_ __dut__.__uuf__._1486_/X __dut__.__uuf__._1480_/X __dut__._2275_/B
+ __dut__.__uuf__._1491_/X __dut__.__uuf__._1493_/X VGND VGND VPWR VPWR __dut__._2274_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2115_ VGND VGND VPWR VPWR __dut__.__uuf__._2115_/HI tie[122] sky130_fd_sc_hd__conb_1
XFILLER_130_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2046_ VGND VGND VPWR VPWR __dut__.__uuf__._2046_/HI tie[53] sky130_fd_sc_hd__conb_1
X__dut__._2300_ __dut__._2300_/A1 __dut__._2300_/A2 __dut__._2299_/X VGND VGND VPWR
+ VPWR __dut__._2300_/X sky130_fd_sc_hd__a21o_4
XFILLER_29_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2231_ __dut__._2325_/A __dut__._2231_/B VGND VGND VPWR VPWR __dut__._2231_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2395__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2162_ __dut__._2172_/A1 __dut__._2162_/A2 __dut__._2161_/X VGND VGND VPWR
+ VPWR __dut__._2162_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2093_ __dut__._2095_/A __dut__._3103_/Q VGND VGND VPWR VPWR __dut__._2093_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_13_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1739__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2995_ __dut__._3093_/CLK __dut__._2995_/D __dut__._2623_/Y VGND VGND VPWR
+ VPWR __dut__._2995_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1946_ __dut__._2172_/A1 tie[125] __dut__._1945_/X VGND VGND VPWR VPWR __dut__._3030_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_125_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1877_ __dut__._1881_/A __dut__._2995_/Q VGND VGND VPWR VPWR __dut__._1877_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2429_ __dut__._2429_/A prod[23] VGND VGND VPWR VPWR __dut__._2429_/X sky130_fd_sc_hd__and2_4
XFILLER_149_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1649__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1504__A2 mp[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1440__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1559__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1615_ __dut__.__uuf__._1615_/A VGND VGND VPWR VPWR __dut__.__uuf__._1615_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1800_ __dut__._1830_/A1 tie[52] __dut__._1799_/X VGND VGND VPWR VPWR __dut__._2957_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1546_ __dut__.__uuf__._1528_/X __dut__.__uuf__._1544_/X __dut__._2249_/B
+ __dut__.__uuf__._1533_/X __dut__.__uuf__._1545_/X VGND VGND VPWR VPWR __dut__._2248_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2780_ rst VGND VGND VPWR VPWR __dut__._2780_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1731_ __dut__._2189_/A __dut__._2922_/Q VGND VGND VPWR VPWR __dut__._1731_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1477_ __dut__._1568_/X __dut__.__uuf__._1465_/X __dut__._2283_/B
+ __dut__.__uuf__._1470_/X VGND VGND VPWR VPWR __dut__.__uuf__._1477_/X sky130_fd_sc_hd__o22a_4
X__dut__._1662_ __dut__._2488_/A1 prod[48] __dut__._1661_/X VGND VGND VPWR VPWR __dut__._2888_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_103_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1593_ __dut__._1593_/A __dut__._2863_/Q VGND VGND VPWR VPWR __dut__._1593_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._2029_ VGND VGND VPWR VPWR __dut__.__uuf__._2029_/HI tie[36] sky130_fd_sc_hd__conb_1
XFILLER_45_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2214_ __dut__._2220_/A1 __dut__._2214_/A2 __dut__._2213_/X VGND VGND VPWR
+ VPWR __dut__._2214_/X sky130_fd_sc_hd__a21o_4
XFILLER_60_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2145_ __dut__._2207_/A __dut__._2145_/B VGND VGND VPWR VPWR __dut__._2145_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_25_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2076_ __dut__._2076_/A1 prod[20] __dut__._2075_/X VGND VGND VPWR VPWR __dut__._3095_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_71_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1469__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2978_ __dut__._3079_/CLK __dut__._2978_/D __dut__._2640_/Y VGND VGND VPWR
+ VPWR __dut__._2978_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1929_ __dut__._2207_/A __dut__._3021_/Q VGND VGND VPWR VPWR __dut__._1929_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_136_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1670__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_112_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2763__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_281 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2141_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_270 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2253_/A sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1379__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_292 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2385_/A sky130_fd_sc_hd__buf_2
XFILLER_145_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1400_ __dut__.__uuf__._1397_/Y __dut__.__uuf__._1398_/X __dut__.__uuf__._1399_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1400_/X sky130_fd_sc_hd__o21a_4
XFILLER_144_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1331_ __dut__.__uuf__._1335_/A VGND VGND VPWR VPWR __dut__.__uuf__._1331_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_116_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1262_ __dut__.__uuf__._1446_/A VGND VGND VPWR VPWR __dut__.__uuf__._1533_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_59_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1193_ __dut__.__uuf__._1192_/X __dut__.__uuf__._1189_/X prod[8]
+ prod[9] __dut__.__uuf__._1185_/X VGND VGND VPWR VPWR __dut__._2398_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._2003__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2673__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._2275__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2901_ __dut__._3109_/CLK __dut__._2901_/D __dut__._2717_/Y VGND VGND VPWR
+ VPWR __dut__._2901_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2832_ clkbuf_5_3_0_tck/X __dut__._2832_/D __dut__._2786_/Y VGND VGND VPWR
+ VPWR __dut__._2832_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2763_ rst VGND VGND VPWR VPWR __dut__._2763_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1529_ __dut__.__uuf__._1550_/A VGND VGND VPWR VPWR __dut__.__uuf__._1529_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_151_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1714_ __dut__._1714_/A1 tie[9] __dut__._1713_/X VGND VGND VPWR VPWR __dut__._2914_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2694_ rst VGND VGND VPWR VPWR __dut__._2694_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_98_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1645_ __dut__._2491_/A __dut__._2879_/Q VGND VGND VPWR VPWR __dut__._1645_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1576_ __dut__._1374_/Y mp[23] __dut__._1575_/X VGND VGND VPWR VPWR __dut__._1576_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_73_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1652__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2583__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2128_ __dut__._2128_/A1 __dut__._2128_/A2 __dut__._2127_/X VGND VGND VPWR
+ VPWR __dut__._2128_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1404__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2059_ __dut__._2407_/A __dut__._3086_/Q VGND VGND VPWR VPWR __dut__._2059_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1927__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._3018__CLK clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2758__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__.__uuf__._1294__A __dut__.__uuf__._1294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1880_ __dut__.__uuf__._1923_/A __dut__.__uuf__._1880_/B __dut__.__uuf__._1880_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1881_/A sky130_fd_sc_hd__or3_4
XFILLER_20_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1837__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2363_ __dut__.__uuf__._2364_/CLK __dut__._2506_/X __dut__.__uuf__._1042_/A
+ VGND VGND VPWR VPWR prod[62] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1469__A __dut__.__uuf__._1533_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1314_ __dut__.__uuf__._1335_/A VGND VGND VPWR VPWR __dut__.__uuf__._1314_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_99_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0_tck clkbuf_3_7_0_tck/A VGND VGND VPWR VPWR clkbuf_3_6_0_tck/X sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2294_ __dut__.__uuf__._2307_/CLK __dut__._2368_/X __dut__.__uuf__._1254_/X
+ VGND VGND VPWR VPWR __dut__._2369_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1245_ __dut__._2375_/B __dut__.__uuf__._1245_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1245_/X sky130_fd_sc_hd__or2_4
XFILLER_143_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2668__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1430_ __dut__._1430_/A1 __dut__._1428_/X __dut__._1429_/X VGND VGND VPWR
+ VPWR __dut__._2823_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1176_ __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR __dut__.__uuf__._1463_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3100_ __dut__._3102_/CLK __dut__._3100_/D __dut__._2518_/Y VGND VGND VPWR
+ VPWR __dut__._3100_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._3031_ clkbuf_5_1_0_tck/X __dut__._3031_/D __dut__._2587_/Y VGND VGND VPWR
+ VPWR __dut__._3031_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_240_ _297_/Q _306_/Q VGND VGND VPWR VPWR _240_/X sky130_fd_sc_hd__or2_4
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_171_ _279_/Q _173_/B VGND VGND VPWR VPWR _278_/D sky130_fd_sc_hd__and2_4
XFILLER_50_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_13_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2815_ __dut__._2509_/B __dut__._2815_/D __dut__._2803_/Y VGND VGND VPWR
+ VPWR __dut__._2815_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1747__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2746_ rst VGND VGND VPWR VPWR __dut__._2746_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2677_ rst VGND VGND VPWR VPWR __dut__._2677_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1628_ __dut__._1374_/Y mc[8] __dut__._1627_/X VGND VGND VPWR VPWR __dut__._1628_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2578__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1559_ __dut__._2509_/A __dut__._2856_/Q VGND VGND VPWR VPWR __dut__._1559_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2050__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1657__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_277_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1030_ __dut__.__uuf__._1992_/A VGND VGND VPWR VPWR __dut__.__uuf__._1042_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_84_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__313__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1616__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1932_ __dut__.__uuf__._1932_/A VGND VGND VPWR VPWR __dut__.__uuf__._1934_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1863_ __dut__.__uuf__._1863_/A VGND VGND VPWR VPWR __dut__.__uuf__._1863_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_149_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1794_ __dut__.__uuf__._1794_/A VGND VGND VPWR VPWR __dut__._2164_/A2
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._1987__B1 __dut__.__uuf__._1023_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1567__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2600_ rst VGND VGND VPWR VPWR __dut__._2600_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2346_ __dut__.__uuf__._2353_/CLK __dut__._2472_/X __dut__.__uuf__._1081_/X
+ VGND VGND VPWR VPWR prod[45] sky130_fd_sc_hd__dfrtp_4
XFILLER_120_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2531_ rst VGND VGND VPWR VPWR __dut__._2531_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2277_ __dut__.__uuf__._2278_/CLK __dut__._2334_/X __dut__.__uuf__._1345_/X
+ VGND VGND VPWR VPWR __dut__._2335_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2462_ __dut__._2488_/A1 __dut__._2462_/A2 __dut__._2461_/X VGND VGND VPWR
+ VPWR __dut__._2462_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1228_ __dut__.__uuf__._1441_/A VGND VGND VPWR VPWR __dut__.__uuf__._1292_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_101_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1413_ __dut__._2189_/A __dut__._2818_/Q VGND VGND VPWR VPWR __dut__._1413_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_47_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1159_ __dut__.__uuf__._1173_/A VGND VGND VPWR VPWR __dut__.__uuf__._1159_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2393_ __dut__._2407_/A prod[5] VGND VGND VPWR VPWR __dut__._2393_/X sky130_fd_sc_hd__and2_4
XFILLER_103_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._3014_ __dut__._3059_/CLK __dut__._3014_/D __dut__._2604_/Y VGND VGND VPWR
+ VPWR __dut__._3014_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_223_ _304_/Q _225_/B VGND VGND VPWR VPWR _297_/D sky130_fd_sc_hd__and2_4
XFILLER_156_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_154_ _238_/A _311_/Q _154_/C _242_/A VGND VGND VPWR VPWR _193_/B sky130_fd_sc_hd__or4_4
XFILLER_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2729_ rst VGND VGND VPWR VPWR __dut__._2729_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__274__CLK _274_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2101__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2771__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1387__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2200_ __dut__.__uuf__._2230_/CLK __dut__._2180_/X __dut__.__uuf__._1601_/X
+ VGND VGND VPWR VPWR __dut__._2181_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_1_0_0___dut__.__uuf__.__clk_source___A clkbuf_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2131_ VGND VGND VPWR VPWR __dut__.__uuf__._2131_/HI tie[138] sky130_fd_sc_hd__conb_1
XFILLER_102_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2062_ VGND VGND VPWR VPWR __dut__.__uuf__._2062_/HI tie[69] sky130_fd_sc_hd__conb_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1013_ __dut__.__uuf__._1226_/A __dut__._2379_/B __dut__._2377_/B
+ __dut__._2375_/B VGND VGND VPWR VPWR __dut__.__uuf__._1014_/D sky130_fd_sc_hd__or4_4
XFILLER_29_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2011__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1915_ __dut__._1440_/X VGND VGND VPWR VPWR __dut__.__uuf__._1919_/B
+ sky130_fd_sc_hd__inv_2
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1846_ __dut__.__uuf__._1813_/X __dut__.__uuf__._1844_/B __dut__.__uuf__._1844_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1847_/C sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._2681__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._1777_ __dut__._2159_/B __dut__._2165_/B VGND VGND VPWR VPWR __dut__.__uuf__._1778_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_137_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1962_ __dut__._2004_/A1 tie[133] __dut__._1961_/X VGND VGND VPWR VPWR __dut__._3038_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1893_ __dut__._2507_/A __dut__._3003_/Q VGND VGND VPWR VPWR __dut__._1893_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_133_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2329_ __dut__.__uuf__._2353_/CLK __dut__._2438_/X __dut__.__uuf__._1131_/X
+ VGND VGND VPWR VPWR prod[28] sky130_fd_sc_hd__dfrtp_4
XFILLER_58_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2873__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2514_ rst VGND VGND VPWR VPWR __dut__._2514_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_80_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2445_ __dut__._2507_/A prod[31] VGND VGND VPWR VPWR __dut__._2445_/X sky130_fd_sc_hd__and2_4
XFILLER_74_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2376_ __dut__._2376_/A1 __dut__._2376_/A2 __dut__._2375_/X VGND VGND VPWR
+ VPWR __dut__._2376_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2209__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2591__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_206_ _206_/A _250_/Q _249_/Q VGND VGND VPWR VPWR _211_/A sky130_fd_sc_hd__or3_4
XFILLER_156_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_137_ _311_/Q VGND VGND VPWR VPWR _238_/B sky130_fd_sc_hd__inv_2
XFILLER_99_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1935__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2492__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_142_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2766__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1700_ __dut__._2131_/B __dut__._2137_/B __dut__.__uuf__._1699_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1701_/C sky130_fd_sc_hd__o21ai_4
X__dut__.__uuf__._1631_ __dut__.__uuf__._1633_/A VGND VGND VPWR VPWR __dut__.__uuf__._1631_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_119_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1562_ __dut__.__uuf__._1562_/A VGND VGND VPWR VPWR __dut__.__uuf__._1562_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1493_ __dut__._1556_/X __dut__.__uuf__._1487_/X __dut__._2277_/B
+ __dut__.__uuf__._1492_/X VGND VGND VPWR VPWR __dut__.__uuf__._1493_/X sky130_fd_sc_hd__o22a_4
XFILLER_115_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2114_ VGND VGND VPWR VPWR __dut__.__uuf__._2114_/HI tie[121] sky130_fd_sc_hd__conb_1
XFILLER_97_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2045_ VGND VGND VPWR VPWR __dut__.__uuf__._2045_/HI tie[52] sky130_fd_sc_hd__conb_1
X__dut__._2230_ __dut__._2230_/A1 __dut__._2230_/A2 __dut__._2229_/X VGND VGND VPWR
+ VPWR __dut__._2230_/X sky130_fd_sc_hd__a21o_4
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2676__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2395__B prod[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2161_ __dut__._2207_/A __dut__._2161_/B VGND VGND VPWR VPWR __dut__._2161_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2092_ __dut__._2092_/A1 prod[28] __dut__._2091_/X VGND VGND VPWR VPWR __dut__._3103_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_100_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1829_ __dut__.__uuf__._1821_/A __dut__.__uuf__._1826_/B __dut__.__uuf__._1828_/X
+ VGND VGND VPWR VPWR __dut__._2174_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_40_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2994_ __dut__._3093_/CLK __dut__._2994_/D __dut__._2624_/Y VGND VGND VPWR
+ VPWR __dut__._2994_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1945_ __dut__._2207_/A __dut__._3029_/Q VGND VGND VPWR VPWR __dut__._1945_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_118_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1876_ __dut__._1876_/A1 tie[90] __dut__._1875_/X VGND VGND VPWR VPWR __dut__._2995_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1755__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3051__CLK __dut__._3059_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2474__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2428_ __dut__._2428_/A1 __dut__._2428_/A2 __dut__._2427_/X VGND VGND VPWR
+ VPWR __dut__._2428_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2181__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2586__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2359_ __dut__._2407_/A __dut__._2359_/B VGND VGND VPWR VPWR __dut__._2359_/X
+ sky130_fd_sc_hd__and2_4
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1850__A __dut__.__uuf__._1904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1665__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_23_0_tck clkbuf_5_23_0_tck/A VGND VGND VPWR VPWR _306_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1440__A2 mc[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1614_ __dut__.__uuf__._1615_/A VGND VGND VPWR VPWR __dut__.__uuf__._1614_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1545_ __dut__._1496_/X __dut__.__uuf__._1529_/X __dut__._2251_/B
+ __dut__.__uuf__._1534_/X VGND VGND VPWR VPWR __dut__.__uuf__._1545_/X sky130_fd_sc_hd__o22a_4
X__dut__._1730_ __dut__._1760_/A1 tie[17] __dut__._1729_/X VGND VGND VPWR VPWR __dut__._2922_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_104_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1575__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1476_ __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR __dut__.__uuf__._1476_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_115_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1661_ __dut__._2491_/A __dut__._2887_/Q VGND VGND VPWR VPWR __dut__._1661_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_39_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1592_ __dut__._1374_/Y mp[27] __dut__._1591_/X VGND VGND VPWR VPWR __dut__._1592_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2028_ VGND VGND VPWR VPWR __dut__.__uuf__._2028_/HI tie[35] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2456__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2213_ __dut__._2507_/A __dut__._2213_/B VGND VGND VPWR VPWR __dut__._2213_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_60_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2144_ __dut__._2144_/A1 __dut__._2144_/A2 __dut__._2143_/X VGND VGND VPWR
+ VPWR __dut__._2144_/X sky130_fd_sc_hd__a21o_4
XFILLER_111_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_43_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2075_ __dut__._2507_/A __dut__._3094_/Q VGND VGND VPWR VPWR __dut__._2075_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_139_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2977_ __dut__._3079_/CLK __dut__._2977_/D __dut__._2641_/Y VGND VGND VPWR
+ VPWR __dut__._2977_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1928_ __dut__._1928_/A1 tie[116] __dut__._1927_/X VGND VGND VPWR VPWR __dut__._3021_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_141_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1859_ __dut__._1881_/A __dut__._2986_/Q VGND VGND VPWR VPWR __dut__._1859_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1554__B2 __dut__.__uuf__._1294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_105_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_271 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2251_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_260 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2269_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_282 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2207_/A sky130_fd_sc_hd__buf_8
XANTENNA___dut__._3097__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_293 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2389_/A sky130_fd_sc_hd__buf_2
XFILLER_145_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1330_ __dut__.__uuf__._1327_/X __dut__.__uuf__._1329_/X __dut__._2343_/B
+ __dut__.__uuf__._1327_/X VGND VGND VPWR VPWR __dut__._2342_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1395__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1261_ __dut__.__uuf__._1921_/A VGND VGND VPWR VPWR __dut__.__uuf__._1261_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1192_ __dut__.__uuf__._1463_/A VGND VGND VPWR VPWR __dut__.__uuf__._1192_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_140_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2934__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._2900_ _306_/CLK __dut__._2900_/D __dut__._2718_/Y VGND VGND VPWR VPWR __dut__._2900_/Q
+ sky130_fd_sc_hd__dfrtp_4
X__dut__._2831_ __dut__._2836_/CLK __dut__._2831_/D __dut__._2787_/Y VGND VGND VPWR
+ VPWR __dut__._2831_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2762_ rst VGND VGND VPWR VPWR __dut__._2762_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1528_ __dut__.__uuf__._1549_/A VGND VGND VPWR VPWR __dut__.__uuf__._1528_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2693_ rst VGND VGND VPWR VPWR __dut__._2693_/Y sky130_fd_sc_hd__inv_2
X__dut__._1713_ __dut__._2189_/A __dut__._2913_/Q VGND VGND VPWR VPWR __dut__._1713_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1459_ __dut__._1584_/X __dut__.__uuf__._1442_/X __dut__._2291_/B
+ __dut__.__uuf__._1448_/X VGND VGND VPWR VPWR __dut__.__uuf__._1459_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1644_ __dut__._2502_/A1 prod[39] __dut__._1643_/X VGND VGND VPWR VPWR __dut__._2879_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_103_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1575_ __dut__._2509_/A __dut__._2860_/Q VGND VGND VPWR VPWR __dut__._1575_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2127_ __dut__._2141_/A __dut__._2127_/B VGND VGND VPWR VPWR __dut__._2127_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1404__A2 mc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2058_ __dut__._2412_/A1 prod[11] __dut__._2057_/X VGND VGND VPWR VPWR __dut__._3086_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_41_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1943__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_222_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2774__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2362_ __dut__.__uuf__._2364_/CLK __dut__._2504_/X __dut__.__uuf__._1032_/X
+ VGND VGND VPWR VPWR prod[61] sky130_fd_sc_hd__dfrtp_4
XFILLER_105_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2293_ __dut__.__uuf__._2293_/CLK __dut__._2366_/X __dut__.__uuf__._1258_/X
+ VGND VGND VPWR VPWR __dut__._2367_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1313_ __dut__.__uuf__._1340_/A VGND VGND VPWR VPWR __dut__.__uuf__._1335_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1244_ __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR __dut__.__uuf__._1244_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_141_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1175_ __dut__.__uuf__._1175_/A VGND VGND VPWR VPWR __dut__.__uuf__._1175_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3030_ clkbuf_5_1_0_tck/X __dut__._3030_/D __dut__._2588_/Y VGND VGND VPWR
+ VPWR __dut__._3030_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2684__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1049__A3 prod[56] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_tck_A tck VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_170_ _280_/Q _172_/B VGND VGND VPWR VPWR _279_/D sky130_fd_sc_hd__or2_4
XFILLER_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2814_ __dut__._2509_/B __dut__._2814_/D __dut__._2804_/Y VGND VGND VPWR
+ VPWR __dut__._2814_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2745_ rst VGND VGND VPWR VPWR __dut__._2745_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2676_ rst VGND VGND VPWR VPWR __dut__._2676_/Y sky130_fd_sc_hd__inv_2
X__dut__._1627_ __dut__._2509_/A __dut__._2873_/Q VGND VGND VPWR VPWR __dut__._1627_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1558_ __dut__._1562_/A1 __dut__._1556_/X __dut__._1557_/X VGND VGND VPWR
+ VPWR __dut__._2855_/D sky130_fd_sc_hd__a21o_4
XFILLER_18_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1489_ __dut__._1493_/A __dut__._2837_/Q VGND VGND VPWR VPWR __dut__._1489_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_93_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2594__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2050__A2 prod[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_299_ _313_/CLK _299_/D trst VGND VGND VPWR VPWR _299_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_127_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2769__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_172_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1673__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2265__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1616__A2 start VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1931_ __dut__.__uuf__._1952_/A __dut__.__uuf__._1931_/B __dut__.__uuf__._1931_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1932_/A sky130_fd_sc_hd__or3_4
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1862_ __dut__._2191_/B __dut__._2197_/B VGND VGND VPWR VPWR __dut__.__uuf__._1863_/A
+ sky130_fd_sc_hd__and2_4
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2009__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1793_ __dut__.__uuf__._1815_/A __dut__.__uuf__._1793_/B __dut__.__uuf__._1793_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1794_/A sky130_fd_sc_hd__or3_4
XFILLER_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2345_ __dut__.__uuf__._2353_/CLK __dut__._2470_/X __dut__.__uuf__._1084_/X
+ VGND VGND VPWR VPWR prod[44] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1552__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2276_ __dut__.__uuf__._2278_/CLK __dut__._2332_/X __dut__.__uuf__._1351_/X
+ VGND VGND VPWR VPWR __dut__._2333_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2679__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2530_ rst VGND VGND VPWR VPWR __dut__._2530_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1583__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2461_ __dut__._2491_/A prod[39] VGND VGND VPWR VPWR __dut__._2461_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1227_ __dut__._2381_/B __dut__.__uuf__._1227_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1227_/X sky130_fd_sc_hd__or2_4
XFILLER_101_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1412_ __dut__._1374_/Y mc[18] __dut__._1411_/X VGND VGND VPWR VPWR __dut__._1412_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1158_ __dut__.__uuf__._1161_/A VGND VGND VPWR VPWR __dut__.__uuf__._1158_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2392_ __dut__._2412_/A1 __dut__._2392_/A2 __dut__._2391_/X VGND VGND VPWR
+ VPWR __dut__._2392_/X sky130_fd_sc_hd__a21o_4
XFILLER_55_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1089_ __dut__.__uuf__._1088_/X __dut__.__uuf__._1085_/X prod[43]
+ prod[44] __dut__.__uuf__._1082_/X VGND VGND VPWR VPWR __dut__._2468_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_103_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3013_ _271_/CLK __dut__._3013_/D __dut__._2605_/Y VGND VGND VPWR VPWR __dut__._3013_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_70_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._3008__CLK _274_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_222_ _222_/A _297_/Q VGND VGND VPWR VPWR _296_/D sky130_fd_sc_hd__and2_4
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_153_ _314_/Q _313_/Q VGND VGND VPWR VPWR _242_/A sky130_fd_sc_hd__or2_4
XFILLER_136_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2728_ rst VGND VGND VPWR VPWR __dut__._2728_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2589__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2659_ rst VGND VGND VPWR VPWR __dut__._2659_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_tck clkbuf_3_5_0_tck/A VGND VGND VPWR VPWR clkbuf_3_5_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2130_ VGND VGND VPWR VPWR __dut__.__uuf__._2130_/HI tie[137] sky130_fd_sc_hd__conb_1
XFILLER_124_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2061_ VGND VGND VPWR VPWR __dut__.__uuf__._2061_/HI tie[68] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1012_ __dut__._2381_/B VGND VGND VPWR VPWR __dut__.__uuf__._1226_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_96_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1914_ __dut__.__uuf__._1907_/A __dut__.__uuf__._1912_/B __dut__.__uuf__._1882_/X
+ VGND VGND VPWR VPWR __dut__._2206_/A2 sky130_fd_sc_hd__o21a_4
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1845_ __dut__.__uuf__._1845_/A VGND VGND VPWR VPWR __dut__.__uuf__._1847_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_33_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1776_ __dut__._1384_/X VGND VGND VPWR VPWR __dut__.__uuf__._1780_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_137_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1961_ __dut__._2005_/A __dut__._3037_/Q VGND VGND VPWR VPWR __dut__._1961_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1892_ __dut__._2004_/A1 tie[98] __dut__._1891_/X VGND VGND VPWR VPWR __dut__._3003_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_133_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2328_ __dut__.__uuf__._2328_/CLK __dut__._2436_/X __dut__.__uuf__._1135_/X
+ VGND VGND VPWR VPWR prod[27] sky130_fd_sc_hd__dfrtp_4
XFILLER_121_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2259_ __dut__.__uuf__._2293_/CLK __dut__._2298_/X __dut__.__uuf__._1434_/X
+ VGND VGND VPWR VPWR __dut__._2299_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2513_ rst VGND VGND VPWR VPWR __dut__._2513_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2444_ __dut__._2444_/A1 __dut__._2444_/A2 __dut__._2443_/X VGND VGND VPWR
+ VPWR __dut__._2444_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_73_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2375_ __dut__._2407_/A __dut__._2375_/B VGND VGND VPWR VPWR __dut__._2375_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_28_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_205_ _248_/Q VGND VGND VPWR VPWR _206_/A sky130_fd_sc_hd__inv_2
XFILLER_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_136_ _312_/Q _138_/B _135_/X _128_/X VGND VGND VPWR VPWR _312_/D sky130_fd_sc_hd__a211o_4
XFILLER_99_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1516__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_6_0_tck_A clkbuf_3_7_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1951__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_135_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2303__CLK __dut__.__uuf__._2303_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2782__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1630_ __dut__.__uuf__._1633_/A VGND VGND VPWR VPWR __dut__.__uuf__._1630_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1561_ __dut__.__uuf__._1549_/X __dut__.__uuf__._1544_/X __dut__._2241_/B
+ __dut__.__uuf__._1447_/A __dut__.__uuf__._1560_/X VGND VGND VPWR VPWR __dut__._2240_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_119_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1492_ __dut__.__uuf__._1492_/A VGND VGND VPWR VPWR __dut__.__uuf__._1492_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_115_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2113_ VGND VGND VPWR VPWR __dut__.__uuf__._2113_/HI tie[120] sky130_fd_sc_hd__conb_1
XFILLER_69_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2044_ VGND VGND VPWR VPWR __dut__.__uuf__._2044_/HI tie[51] sky130_fd_sc_hd__conb_1
XFILLER_29_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2160_ __dut__._2172_/A1 __dut__._2160_/A2 __dut__._2159_/X VGND VGND VPWR
+ VPWR __dut__._2160_/X sky130_fd_sc_hd__a21o_4
XANTENNA__241__A1 tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2091_ __dut__._2095_/A __dut__._3102_/Q VGND VGND VPWR VPWR __dut__._2091_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_25_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1994__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2692__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1828_ __dut__.__uuf__._1828_/A VGND VGND VPWR VPWR __dut__.__uuf__._1828_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_40_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2993_ __dut__._3093_/CLK __dut__._2993_/D __dut__._2625_/Y VGND VGND VPWR
+ VPWR __dut__._2993_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1759_ __dut__.__uuf__._1982_/A VGND VGND VPWR VPWR __dut__.__uuf__._1759_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_153_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1944_ __dut__._2172_/A1 tie[124] __dut__._1943_/X VGND VGND VPWR VPWR __dut__._3029_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_109_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1875_ __dut__._1881_/A __dut__._2994_/Q VGND VGND VPWR VPWR __dut__._1875_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2990__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_7_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2427_ __dut__._2427_/A prod[22] VGND VGND VPWR VPWR __dut__._2427_/X sky130_fd_sc_hd__and2_4
XFILLER_85_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2358_ __dut__._2368_/A1 __dut__._2358_/A2 __dut__._2357_/X VGND VGND VPWR
+ VPWR __dut__._2358_/X sky130_fd_sc_hd__a21o_4
X__dut__._2289_ __dut__._2303_/A __dut__._2289_/B VGND VGND VPWR VPWR __dut__._2289_/X
+ sky130_fd_sc_hd__and2_4
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2107__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0___dut__.__uuf__.__clk_source__ clkbuf_4_9_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2328_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_144_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2162__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2777__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_252_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__287__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0___dut__.__uuf__.__clk_source__ clkbuf_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR clkbuf_2_1_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1976__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2017__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1613_ __dut__.__uuf__._1615_/A VGND VGND VPWR VPWR __dut__.__uuf__._1613_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1544_ __dut__.__uuf__._1563_/A VGND VGND VPWR VPWR __dut__.__uuf__._1544_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1475_ __dut__.__uuf__._1463_/X __dut__.__uuf__._1458_/X __dut__._2283_/B
+ __dut__.__uuf__._1469_/X __dut__.__uuf__._1474_/X VGND VGND VPWR VPWR __dut__._2282_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_89_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1660_ __dut__._2488_/A1 prod[47] __dut__._1659_/X VGND VGND VPWR VPWR __dut__._2887_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1900__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1591_ __dut__._2509_/A __dut__._2864_/Q VGND VGND VPWR VPWR __dut__._1591_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2027_ VGND VGND VPWR VPWR __dut__.__uuf__._2027_/HI tie[34] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2687__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1591__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2212_ __dut__._2212_/A1 __dut__._2212_/A2 __dut__._2211_/X VGND VGND VPWR
+ VPWR __dut__._2212_/X sky130_fd_sc_hd__a21o_4
XFILLER_38_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2143_ __dut__._2207_/A __dut__._2143_/B VGND VGND VPWR VPWR __dut__._2143_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_111_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_36_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2074_ __dut__._2074_/A1 prod[19] __dut__._2073_/X VGND VGND VPWR VPWR __dut__._3094_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2392__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2976_ __dut__._3079_/CLK __dut__._2976_/D __dut__._2642_/Y VGND VGND VPWR
+ VPWR __dut__._2976_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1927_ __dut__._2207_/A __dut__._3020_/Q VGND VGND VPWR VPWR __dut__._1927_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_107_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1858_ __dut__._1864_/A1 tie[81] __dut__._1857_/X VGND VGND VPWR VPWR __dut__._2986_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_136_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1789_ __dut__._1797_/A __dut__._2951_/Q VGND VGND VPWR VPWR __dut__._1789_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2597__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2886__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpsn_inst_psn_buff_250 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1593_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_272 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2249_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_261 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2267_/A sky130_fd_sc_hd__buf_2
XFILLER_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_294 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2415_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_283 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2245_/A sky130_fd_sc_hd__buf_2
XFILLER_117_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__307__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1260_ __dut__.__uuf__._1703_/A VGND VGND VPWR VPWR __dut__.__uuf__._1921_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1191_ __dut__.__uuf__._1191_/A VGND VGND VPWR VPWR __dut__.__uuf__._1191_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_140_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_3_0_tck_A clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1233__A1 __dut__.__uuf__._1214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2830_ __dut__._2836_/CLK __dut__._2830_/D __dut__._2788_/Y VGND VGND VPWR
+ VPWR __dut__._2830_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2171__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1527_ __dut__.__uuf__._1543_/A VGND VGND VPWR VPWR __dut__.__uuf__._1527_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2761_ rst VGND VGND VPWR VPWR __dut__._2761_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2692_ rst VGND VGND VPWR VPWR __dut__._2692_/Y sky130_fd_sc_hd__inv_2
X__dut__._1712_ __dut__._1714_/A1 tie[8] __dut__._1711_/X VGND VGND VPWR VPWR __dut__._2913_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1458_ __dut__.__uuf__._1480_/A VGND VGND VPWR VPWR __dut__.__uuf__._1458_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1643_ __dut__._2457_/A __dut__._2878_/Q VGND VGND VPWR VPWR __dut__._1643_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1389_ __dut__.__uuf__._1414_/A VGND VGND VPWR VPWR __dut__.__uuf__._1389_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_106_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1574_ __dut__._1780_/A1 __dut__._1572_/X __dut__._1573_/X VGND VGND VPWR
+ VPWR __dut__._2859_/D sky130_fd_sc_hd__a21o_4
XFILLER_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2126_ __dut__._2126_/A1 __dut__._2126_/A2 __dut__._2125_/X VGND VGND VPWR
+ VPWR __dut__._2126_/X sky130_fd_sc_hd__a21o_4
XANTENNA_clkbuf_4_5_0_tck_A clkbuf_4_5_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2057_ __dut__._2407_/A __dut__._3085_/Q VGND VGND VPWR VPWR __dut__._2057_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_5_22_0_tck clkbuf_5_23_0_tck/A VGND VGND VPWR VPWR __dut__._3109_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_142_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2959_ __dut__._2985_/CLK __dut__._2959_/D __dut__._2659_/Y VGND VGND VPWR
+ VPWR __dut__._2959_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._3064__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_215_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2790__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1215__A1 __dut__.__uuf__._1206_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2194__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2356__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2901__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2361_ __dut__.__uuf__._2364_/CLK __dut__._2502_/X __dut__.__uuf__._1034_/X
+ VGND VGND VPWR VPWR prod[60] sky130_fd_sc_hd__dfrtp_4
XFILLER_145_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2292_ __dut__.__uuf__._2293_/CLK __dut__._2364_/X __dut__.__uuf__._1265_/X
+ VGND VGND VPWR VPWR __dut__._2365_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1312_ __dut__.__uuf__._1300_/X __dut__.__uuf__._1310_/X __dut__._2349_/B
+ __dut__.__uuf__._1311_/X VGND VGND VPWR VPWR __dut__._2348_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1243_ __dut__.__uuf__._1254_/A VGND VGND VPWR VPWR __dut__.__uuf__._1243_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_99_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1174_ __dut__.__uuf__._1162_/X __dut__.__uuf__._1173_/X prod[14]
+ prod[15] __dut__.__uuf__._1170_/X VGND VGND VPWR VPWR __dut__._2410_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_100_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2813_ clkbuf_5_9_0_tck/X __dut__._2813_/D __dut__._2805_/Y VGND VGND VPWR
+ VPWR __dut__._2813_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2205__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2744_ rst VGND VGND VPWR VPWR __dut__._2744_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2675_ rst VGND VGND VPWR VPWR __dut__._2675_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1626_ __dut__._1626_/A1 __dut__._1624_/X __dut__._1625_/X VGND VGND VPWR
+ VPWR __dut__._2872_/D sky130_fd_sc_hd__a21o_4
XFILLER_77_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1557_ __dut__._1557_/A __dut__._2853_/Q VGND VGND VPWR VPWR __dut__._1557_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_100_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3087__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1693__A1 __dut__.__uuf__._1261_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1488_ __dut__._1374_/Y mp[3] __dut__._1487_/X VGND VGND VPWR VPWR __dut__._1488_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_18_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2109_ __dut__._2325_/A __dut__._2109_/B VGND VGND VPWR VPWR __dut__._2109_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2924__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._3089_ __dut__._3093_/CLK __dut__._3089_/D __dut__._2529_/Y VGND VGND VPWR
+ VPWR __dut__._3089_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2338__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_298_ _313_/CLK _298_/D trst VGND VGND VPWR VPWR _298_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2115__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2510__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_165_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2785__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1930_ __dut__._2215_/B __dut__._2221_/B __dut__.__uuf__._1929_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1931_/C sky130_fd_sc_hd__o21ai_4
X__dut__.__uuf__._1861_ __dut__._1416_/X VGND VGND VPWR VPWR __dut__.__uuf__._1865_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1792_ __dut__.__uuf__._1759_/X __dut__.__uuf__._1790_/B __dut__.__uuf__._1790_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1793_/C sky130_fd_sc_hd__o21a_4
XFILLER_137_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2025__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2344_ __dut__.__uuf__._2353_/CLK __dut__._2468_/X __dut__.__uuf__._1087_/X
+ VGND VGND VPWR VPWR prod[43] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1552__A2 mc[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2275_ __dut__.__uuf__._2278_/CLK __dut__._2330_/X __dut__.__uuf__._1356_/X
+ VGND VGND VPWR VPWR __dut__._2331_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2460_ __dut__._2502_/A1 __dut__._2460_/A2 __dut__._2459_/X VGND VGND VPWR
+ VPWR __dut__._2460_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1226_ __dut__.__uuf__._1226_/A __dut__.__uuf__._1226_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1226_/X sky130_fd_sc_hd__or2_4
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1411_ __dut__._2509_/A __dut__._2819_/Q VGND VGND VPWR VPWR __dut__._1411_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1157_ __dut__.__uuf__._1147_/X __dut__.__uuf__._1144_/X prod[20]
+ prod[21] __dut__.__uuf__._1156_/X VGND VGND VPWR VPWR __dut__._2422_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_101_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_0_0_tck_A clkbuf_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2391_ __dut__._2391_/A prod[4] VGND VGND VPWR VPWR __dut__._2391_/X sky130_fd_sc_hd__and2_4
XFILLER_74_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2695__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1088_ __dut__.__uuf__._1088_/A VGND VGND VPWR VPWR __dut__.__uuf__._1088_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1124__B1 prod[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._3012_ _271_/CLK __dut__._3012_/D __dut__._2606_/Y VGND VGND VPWR VPWR __dut__._3012_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_221_ _292_/Q _220_/A _222_/A VGND VGND VPWR VPWR _295_/D sky130_fd_sc_hd__o21a_4
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_152_ _302_/Q VGND VGND VPWR VPWR _154_/C sky130_fd_sc_hd__inv_2
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2727_ rst VGND VGND VPWR VPWR __dut__._2727_/Y sky130_fd_sc_hd__inv_2
X__dut__._2658_ rst VGND VGND VPWR VPWR __dut__._2658_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1609_ __dut__._1609_/A __dut__._2867_/Q VGND VGND VPWR VPWR __dut__._1609_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_93_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2589_ rst VGND VGND VPWR VPWR __dut__._2589_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0___dut__.__uuf__.__clk_source__ clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_3_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_119_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3102__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1949__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2232__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_282_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2060_ VGND VGND VPWR VPWR __dut__.__uuf__._2060_/HI tie[67] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2499__B prod[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1011_ __dut__._2371_/B VGND VGND VPWR VPWR __dut__.__uuf__._1219_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_13_0_tck_A clkbuf_3_6_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1913_ __dut__.__uuf__._1913_/A VGND VGND VPWR VPWR __dut__._2208_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1844_ __dut__.__uuf__._1844_/A __dut__.__uuf__._1844_/B __dut__.__uuf__._1844_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1845_/A sky130_fd_sc_hd__or3_4
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1775_ __dut__.__uuf__._1767_/A __dut__.__uuf__._1772_/B __dut__.__uuf__._1774_/X
+ VGND VGND VPWR VPWR __dut__._2154_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1960_ __dut__._1960_/A1 tie[132] __dut__._1959_/X VGND VGND VPWR VPWR __dut__._3037_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_137_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1891_ __dut__._1891_/A __dut__._3002_/Q VGND VGND VPWR VPWR __dut__._1891_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_133_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2327_ __dut__.__uuf__._2353_/CLK __dut__._2434_/X __dut__.__uuf__._1137_/X
+ VGND VGND VPWR VPWR prod[26] sky130_fd_sc_hd__dfrtp_4
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2258_ __dut__.__uuf__._2293_/CLK __dut__._2296_/X __dut__.__uuf__._1439_/X
+ VGND VGND VPWR VPWR __dut__._2297_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2512_ rst VGND VGND VPWR VPWR __dut__._2512_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1209_ __dut__.__uuf__._1234_/A VGND VGND VPWR VPWR __dut__.__uuf__._1209_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_75_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2443_ __dut__._2507_/A prod[30] VGND VGND VPWR VPWR __dut__._2443_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._2189_ __dut__.__uuf__._2216_/CLK __dut__._2158_/X __dut__.__uuf__._1615_/X
+ VGND VGND VPWR VPWR __dut__._2159_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2374_ __dut__._2376_/A1 __dut__._2374_/A2 __dut__._2373_/X VGND VGND VPWR
+ VPWR __dut__._2374_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_66_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1112__A3 prod[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_204_ _246_/Q VGND VGND VPWR VPWR _204_/Y sky130_fd_sc_hd__inv_2
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_135_ _308_/Q _231_/A VGND VGND VPWR VPWR _135_/X sky130_fd_sc_hd__and2_4
Xclkbuf_4_15_0_tck clkbuf_3_7_0_tck/X VGND VGND VPWR VPWR clkbuf_5_31_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_99_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1516__A2 mp[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_128_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1452__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1560_ __dut__._1480_/X __dut__.__uuf__._1550_/X __dut__._2243_/B
+ __dut__.__uuf__._1294_/A VGND VGND VPWR VPWR __dut__.__uuf__._1560_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1491_ __dut__.__uuf__._1533_/A VGND VGND VPWR VPWR __dut__.__uuf__._1491_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2112_ VGND VGND VPWR VPWR __dut__.__uuf__._2112_/HI tie[119] sky130_fd_sc_hd__conb_1
XFILLER_69_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2043_ VGND VGND VPWR VPWR __dut__.__uuf__._2043_/HI tie[50] sky130_fd_sc_hd__conb_1
XFILLER_57_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1774__A __dut__.__uuf__._1828_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2090_ __dut__._2488_/A1 prod[27] __dut__._2089_/X VGND VGND VPWR VPWR __dut__._3102_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_25_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1827_ __dut__.__uuf__._1827_/A VGND VGND VPWR VPWR __dut__._2176_/A2
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2278__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_138_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2992_ __dut__._3093_/CLK __dut__._2992_/D __dut__._2626_/Y VGND VGND VPWR
+ VPWR __dut__._2992_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1758_ __dut__.__uuf__._1758_/A VGND VGND VPWR VPWR __dut__.__uuf__._1761_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1689_ __dut__.__uuf__._1689_/A VGND VGND VPWR VPWR __dut__.__uuf__._1689_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1943_ __dut__._2189_/A __dut__._3028_/Q VGND VGND VPWR VPWR __dut__._1943_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_109_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1874_ __dut__._1874_/A1 tie[89] __dut__._1873_/X VGND VGND VPWR VPWR __dut__._2994_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2213__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_tck clkbuf_3_5_0_tck/A VGND VGND VPWR VPWR clkbuf_4_9_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_125_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2426_ __dut__._2426_/A1 __dut__._2426_/A2 __dut__._2425_/X VGND VGND VPWR
+ VPWR __dut__._2426_/X sky130_fd_sc_hd__a21o_4
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1682__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2357_ __dut__._2407_/A __dut__._2357_/B VGND VGND VPWR VPWR __dut__._2357_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2288_ __dut__._2288_/A1 __dut__._2288_/A2 __dut__._2287_/X VGND VGND VPWR
+ VPWR __dut__._2288_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1499__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2123__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_245_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2793__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1612_ __dut__.__uuf__._1615_/A VGND VGND VPWR VPWR __dut__.__uuf__._1612_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1543_ __dut__.__uuf__._1543_/A VGND VGND VPWR VPWR __dut__.__uuf__._1543_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1474_ __dut__._1572_/X __dut__.__uuf__._1465_/X __dut__._2285_/B
+ __dut__.__uuf__._1470_/X VGND VGND VPWR VPWR __dut__.__uuf__._1474_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__._2033__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1590_ __dut__._1780_/A1 __dut__._1588_/X __dut__._1589_/X VGND VGND VPWR
+ VPWR __dut__._2863_/D sky130_fd_sc_hd__a21o_4
XFILLER_39_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2026_ VGND VGND VPWR VPWR __dut__.__uuf__._2026_/HI tie[33] sky130_fd_sc_hd__conb_1
XFILLER_84_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1664__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2211_ __dut__._2507_/A __dut__._2211_/B VGND VGND VPWR VPWR __dut__._2211_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._3014__D __dut__._3014_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2142_ __dut__._2142_/A1 __dut__._2142_/A2 __dut__._2141_/X VGND VGND VPWR
+ VPWR __dut__._2142_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1416__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2073_ __dut__._2073_/A __dut__._3093_/Q VGND VGND VPWR VPWR __dut__._2073_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_25_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_29_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2975_ __dut__._2985_/CLK __dut__._2975_/D __dut__._2643_/Y VGND VGND VPWR
+ VPWR __dut__._2975_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1926_ __dut__._1926_/A1 tie[115] __dut__._1925_/X VGND VGND VPWR VPWR __dut__._3020_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_153_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1857_ __dut__._1881_/A __dut__._2985_/Q VGND VGND VPWR VPWR __dut__._1857_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1788_ __dut__._1788_/A1 tie[46] __dut__._1787_/X VGND VGND VPWR VPWR __dut__._2951_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2409_ __dut__._2415_/A prod[13] VGND VGND VPWR VPWR __dut__._2409_/X sky130_fd_sc_hd__and2_4
XFILLER_90_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_240 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1805_/A sky130_fd_sc_hd__buf_2
XFILLER_31_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_262 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2265_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_251 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1601_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_273 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2247_/A sky130_fd_sc_hd__buf_2
XFILLER_129_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_284 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2197_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_295 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2103_/A sky130_fd_sc_hd__buf_2
XFILLER_144_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1957__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1894__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1190_ __dut__.__uuf__._1177_/X __dut__.__uuf__._1189_/X prod[9]
+ prod[10] __dut__.__uuf__._1185_/X VGND VGND VPWR VPWR __dut__._2400_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._2788__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1646__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1526_ __dut__.__uuf__._1566_/A VGND VGND VPWR VPWR __dut__.__uuf__._1543_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_135_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2760_ rst VGND VGND VPWR VPWR __dut__._2760_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1711_ __dut__._2189_/A __dut__._2912_/Q VGND VGND VPWR VPWR __dut__._1711_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2691_ rst VGND VGND VPWR VPWR __dut__._2691_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1457_ __dut__.__uuf__._1457_/A VGND VGND VPWR VPWR __dut__.__uuf__._1457_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_104_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1388_ __dut__.__uuf__._1387_/Y __dut__.__uuf__._1373_/X __dut__.__uuf__._1374_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1388_/X sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._2698__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1642_ __dut__._2502_/A1 prod[38] __dut__._1641_/X VGND VGND VPWR VPWR __dut__._2878_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_131_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1573_ __dut__._1573_/A __dut__._2858_/Q VGND VGND VPWR VPWR __dut__._1573_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_85_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2009_ VGND VGND VPWR VPWR __dut__.__uuf__._2009_/HI tie[16] sky130_fd_sc_hd__conb_1
XFILLER_18_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__.__uuf__._1962__A __dut__.__uuf__._1982_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2125_ __dut__._2325_/A __dut__._2125_/B VGND VGND VPWR VPWR __dut__._2125_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_13_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2062__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2056_ __dut__._2412_/A1 prod[10] __dut__._2055_/X VGND VGND VPWR VPWR __dut__._3085_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_139_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2958_ __dut__._2958_/CLK __dut__._2958_/D __dut__._2660_/Y VGND VGND VPWR
+ VPWR __dut__._2958_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1909_ __dut__._2005_/A __dut__._3011_/Q VGND VGND VPWR VPWR __dut__._1909_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2889_ __dut__._3102_/CLK __dut__._2889_/D __dut__._2729_/Y VGND VGND VPWR
+ VPWR __dut__._2889_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2853__CLK __dut__._2860_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2401__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1628__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_110_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_208_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2360_ __dut__.__uuf__._2364_/CLK __dut__._2500_/X __dut__.__uuf__._1038_/X
+ VGND VGND VPWR VPWR prod[59] sky130_fd_sc_hd__dfrtp_4
XFILLER_132_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2291_ __dut__.__uuf__._2291_/CLK __dut__._2362_/X __dut__.__uuf__._1270_/X
+ VGND VGND VPWR VPWR __dut__._2363_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1311_ __dut__.__uuf__._1311_/A VGND VGND VPWR VPWR __dut__.__uuf__._1311_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1242_ __dut__.__uuf__._1240_/Y __dut__.__uuf__._1241_/X __dut__.__uuf__._1214_/X
+ __dut__._2377_/B __dut__.__uuf__._1232_/X VGND VGND VPWR VPWR __dut__._2376_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_113_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1173_ __dut__.__uuf__._1173_/A VGND VGND VPWR VPWR __dut__.__uuf__._1173_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2311__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2812_ clkbuf_5_2_0_tck/X __dut__._2812_/D __dut__._2806_/Y VGND VGND VPWR
+ VPWR __dut__._2812_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1509_ __dut__._1536_/X __dut__.__uuf__._1508_/X __dut__._2269_/B
+ __dut__.__uuf__._1492_/X VGND VGND VPWR VPWR __dut__.__uuf__._1509_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__.__uuf__._1022__A __dut__.__uuf__._1464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2743_ rst VGND VGND VPWR VPWR __dut__._2743_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2876__CLK __dut__._3109_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2674_ rst VGND VGND VPWR VPWR __dut__._2674_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1625_ __dut__._2197_/A __dut__._2871_/Q VGND VGND VPWR VPWR __dut__._1625_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_96_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2221__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1556_ __dut__._1374_/Y mp[18] __dut__._1555_/X VGND VGND VPWR VPWR __dut__._1556_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_133_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1487_ __dut__._2509_/A __dut__._2838_/Q VGND VGND VPWR VPWR __dut__._1487_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2108_ __dut__._2376_/A1 __dut__._2108_/A2 __dut__._2107_/X VGND VGND VPWR
+ VPWR __dut__._2108_/X sky130_fd_sc_hd__a21o_4
X__dut__._3088_ __dut__._3106_/CLK __dut__._3088_/D __dut__._2530_/Y VGND VGND VPWR
+ VPWR __dut__._3088_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2039_ __dut__._2039_/A __dut__._3076_/Q VGND VGND VPWR VPWR __dut__._2039_/X
+ sky130_fd_sc_hd__and2_4
X_297_ _306_/CLK _297_/D trst VGND VGND VPWR VPWR _297_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_114_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2510__A2 clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_158_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._3031__CLK clkbuf_5_1_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1860_ __dut__.__uuf__._1853_/A __dut__.__uuf__._1858_/B __dut__.__uuf__._1828_/X
+ VGND VGND VPWR VPWR __dut__._2186_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1436__A2 __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1791_ __dut__.__uuf__._1791_/A VGND VGND VPWR VPWR __dut__.__uuf__._1793_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_149_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2343_ __dut__.__uuf__._2353_/CLK __dut__._2466_/X __dut__.__uuf__._1091_/X
+ VGND VGND VPWR VPWR prod[42] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2274_ __dut__.__uuf__._2278_/CLK __dut__._2328_/X __dut__.__uuf__._1360_/X
+ VGND VGND VPWR VPWR __dut__._2329_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_87_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1225_ __dut__.__uuf__._1227_/B VGND VGND VPWR VPWR __dut__.__uuf__._1226_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1410_ __dut__._1410_/A1 __dut__._1408_/X __dut__._1409_/X VGND VGND VPWR
+ VPWR __dut__._2818_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1156_ __dut__.__uuf__._1200_/A VGND VGND VPWR VPWR __dut__.__uuf__._1156_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2390_ __dut__._2412_/A1 __dut__._2390_/A2 __dut__._2389_/X VGND VGND VPWR
+ VPWR __dut__._2390_/X sky130_fd_sc_hd__a21o_4
XFILLER_86_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1087_ __dut__.__uuf__._1087_/A VGND VGND VPWR VPWR __dut__.__uuf__._1087_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_21_0_tck clkbuf_5_21_0_tck/A VGND VGND VPWR VPWR __dut__._3106_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._3011_ _274_/CLK __dut__._3011_/D __dut__._2607_/Y VGND VGND VPWR VPWR __dut__._3011_/Q
+ sky130_fd_sc_hd__dfrtp_4
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1017__A __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_220_ _220_/A _225_/B VGND VGND VPWR VPWR _294_/D sky130_fd_sc_hd__and2_4
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1989_ __dut__.__uuf__._1989_/A __dut__._2109_/B __dut__.__uuf__._1989_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1990_/A sky130_fd_sc_hd__or3_4
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_151_ _312_/Q VGND VGND VPWR VPWR _238_/A sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_11_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3054__CLK __dut__._3059_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2726_ rst VGND VGND VPWR VPWR __dut__._2726_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2657_ rst VGND VGND VPWR VPWR __dut__._2657_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1608_ __dut__._1374_/Y mp[30] __dut__._1607_/X VGND VGND VPWR VPWR __dut__._1608_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2184__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2588_ rst VGND VGND VPWR VPWR __dut__._2588_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1539_ __dut__._2509_/A __dut__._2851_/Q VGND VGND VPWR VPWR __dut__._1539_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_275_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1010_ __dut__._2107_/B VGND VGND VPWR VPWR __dut__.__uuf__._1989_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_110_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2796__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1912_ __dut__.__uuf__._1923_/A __dut__.__uuf__._1912_/B __dut__.__uuf__._1912_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1913_/A sky130_fd_sc_hd__or3_4
XFILLER_37_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1843_ __dut__._2183_/B __dut__._2189_/B __dut__.__uuf__._1842_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1844_/C sky130_fd_sc_hd__o21ai_4
XFILLER_138_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1774_ __dut__.__uuf__._1828_/A VGND VGND VPWR VPWR __dut__.__uuf__._1774_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1890_ __dut__._2502_/A1 tie[97] __dut__._1889_/X VGND VGND VPWR VPWR __dut__._3002_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_145_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2326_ __dut__.__uuf__._2353_/CLK __dut__._2432_/X __dut__.__uuf__._1139_/X
+ VGND VGND VPWR VPWR prod[25] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2257_ __dut__.__uuf__._2293_/CLK __dut__._2294_/X __dut__.__uuf__._1445_/X
+ VGND VGND VPWR VPWR __dut__._2295_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2511_ rst VGND VGND VPWR VPWR __dut__._2511_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2486__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1208_ __dut__.__uuf__._1208_/A VGND VGND VPWR VPWR __dut__.__uuf__._1234_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2914__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2442_ __dut__._2442_/A1 __dut__._2442_/A2 __dut__._2441_/X VGND VGND VPWR
+ VPWR __dut__._2442_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2188_ __dut__.__uuf__._2216_/CLK __dut__._2156_/X __dut__.__uuf__._1617_/X
+ VGND VGND VPWR VPWR __dut__._2157_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_75_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1139_ __dut__.__uuf__._1146_/A VGND VGND VPWR VPWR __dut__.__uuf__._1139_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2373_ __dut__._2407_/A __dut__._2373_/B VGND VGND VPWR VPWR __dut__._2373_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_28_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_59_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_203_ _203_/A VGND VGND VPWR VPWR _203_/X sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2410__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_134_ _134_/A VGND VGND VPWR VPWR _313_/D sky130_fd_sc_hd__inv_2
XFILLER_137_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1033__B1 prod[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2709_ rst VGND VGND VPWR VPWR __dut__._2709_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1988__B1 __dut__._1987_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1452__A2 mc[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1695__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1490_ __dut__.__uuf__._1501_/A VGND VGND VPWR VPWR __dut__.__uuf__._1490_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_127_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2111_ VGND VGND VPWR VPWR __dut__.__uuf__._2111_/HI tie[118] sky130_fd_sc_hd__conb_1
XFILLER_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2042_ VGND VGND VPWR VPWR __dut__.__uuf__._2042_/HI tie[49] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2468__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1826_ __dut__.__uuf__._1869_/A __dut__.__uuf__._1826_/B __dut__.__uuf__._1826_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1827_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1757_ __dut__.__uuf__._1790_/A __dut__.__uuf__._1757_/B __dut__.__uuf__._1757_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1758_/A sky130_fd_sc_hd__or3_4
X__dut__._2991_ __dut__._3093_/CLK __dut__._2991_/D __dut__._2627_/Y VGND VGND VPWR
+ VPWR __dut__._2991_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1688_ __dut__._2127_/B __dut__._2133_/B VGND VGND VPWR VPWR __dut__.__uuf__._1689_/A
+ sky130_fd_sc_hd__and2_4
X__dut__._1942_ __dut__._1942_/A1 tie[123] __dut__._1941_/X VGND VGND VPWR VPWR __dut__._3028_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1873_ __dut__._1881_/A __dut__._2993_/Q VGND VGND VPWR VPWR __dut__._1873_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_109_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1030__A __dut__.__uuf__._1992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2309_ __dut__.__uuf__._2334_/CLK __dut__._2398_/X __dut__.__uuf__._1191_/X
+ VGND VGND VPWR VPWR prod[8] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2425_ __dut__._2507_/A prod[21] VGND VGND VPWR VPWR __dut__._2425_/X sky130_fd_sc_hd__and2_4
XFILLER_75_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1682__A2 prod[58] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2356_ __dut__._2368_/A1 __dut__._2356_/A2 __dut__._2355_/X VGND VGND VPWR
+ VPWR __dut__._2356_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2287_ __dut__._2303_/A __dut__._2287_/B VGND VGND VPWR VPWR __dut__._2287_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1557__B2 __dut__.__uuf__._1294_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_140_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_238_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1611_ __dut__.__uuf__._1615_/A VGND VGND VPWR VPWR __dut__.__uuf__._1611_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1542_ __dut__.__uuf__._1528_/X __dut__.__uuf__._1523_/X __dut__._2251_/B
+ __dut__.__uuf__._1533_/X __dut__.__uuf__._1541_/X VGND VGND VPWR VPWR __dut__._2250_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1473_ __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR __dut__.__uuf__._1473_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_116_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2025_ VGND VGND VPWR VPWR __dut__.__uuf__._2025_/HI tie[32] sky130_fd_sc_hd__conb_1
X__dut__._2210_ __dut__._2212_/A1 __dut__._2210_/A2 __dut__._2209_/X VGND VGND VPWR
+ VPWR __dut__._2210_/X sky130_fd_sc_hd__a21o_4
XFILLER_57_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2141_ __dut__._2141_/A __dut__._2141_/B VGND VGND VPWR VPWR __dut__._2141_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1416__A2 mc[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_14_0_tck clkbuf_3_7_0_tck/X VGND VGND VPWR VPWR clkbuf_5_29_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2072_ __dut__._2422_/A1 prod[18] __dut__._2071_/X VGND VGND VPWR VPWR __dut__._3093_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_111_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1025__A __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1809_ __dut__.__uuf__._1809_/A VGND VGND VPWR VPWR __dut__.__uuf__._1809_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_154_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2974_ __dut__._2985_/CLK __dut__._2974_/D __dut__._2644_/Y VGND VGND VPWR
+ VPWR __dut__._2974_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1925_ __dut__._2207_/A __dut__._3019_/Q VGND VGND VPWR VPWR __dut__._1925_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_138_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1856_ __dut__._1864_/A1 tie[80] __dut__._1855_/X VGND VGND VPWR VPWR __dut__._2985_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1787_ __dut__._1787_/A __dut__._2950_/Q VGND VGND VPWR VPWR __dut__._1787_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2408_ __dut__._2412_/A1 __dut__._2408_/A2 __dut__._2407_/X VGND VGND VPWR
+ VPWR __dut__._2408_/X sky130_fd_sc_hd__a21o_4
XFILLER_29_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0___dut__.__uuf__.__clk_source___A clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2339_ __dut__._2407_/A __dut__._2339_/B VGND VGND VPWR VPWR __dut__._2339_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_230 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2035_/A sky130_fd_sc_hd__buf_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_241 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1807_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_263 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1493_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_252 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1605_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_285 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1557_/A sky130_fd_sc_hd__buf_2
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_274 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1429_/A sky130_fd_sc_hd__buf_2
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_296 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1689_/A sky130_fd_sc_hd__buf_2
XFILLER_117_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1973__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2268__CLK __dut__.__uuf__._2278_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2309__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_tck clkbuf_3_3_0_tck/A VGND VGND VPWR VPWR clkbuf_4_7_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_136_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1525_ __dut__.__uuf__._1507_/X __dut__.__uuf__._1523_/X __dut__._2259_/B
+ __dut__.__uuf__._1512_/X __dut__.__uuf__._1524_/X VGND VGND VPWR VPWR __dut__._2258_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_135_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1710_ __dut__._1714_/A1 tie[7] __dut__._1709_/X VGND VGND VPWR VPWR __dut__._2912_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2690_ rst VGND VGND VPWR VPWR __dut__._2690_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1456_ __dut__.__uuf__._1440_/X __dut__.__uuf__._1435_/X __dut__._2291_/B
+ __dut__.__uuf__._1447_/X __dut__.__uuf__._1455_/X VGND VGND VPWR VPWR __dut__._2290_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_150_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1387_ __dut__._2321_/B VGND VGND VPWR VPWR __dut__.__uuf__._1387_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1641_ __dut__._2457_/A __dut__._2877_/Q VGND VGND VPWR VPWR __dut__._1641_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_131_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1572_ __dut__._1374_/Y mp[22] __dut__._1571_/X VGND VGND VPWR VPWR __dut__._1572_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_85_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2008_ VGND VGND VPWR VPWR __dut__.__uuf__._2008_/HI tie[15] sky130_fd_sc_hd__conb_1
XFILLER_122_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2124_ __dut__._2332_/A1 __dut__._2124_/A2 __dut__._2123_/X VGND VGND VPWR
+ VPWR __dut__._2124_/X sky130_fd_sc_hd__a21o_4
XFILLER_82_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2219__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_41_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2055_ __dut__._2407_/A __dut__._3084_/Q VGND VGND VPWR VPWR __dut__._2055_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_139_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2957_ __dut__._2958_/CLK __dut__._2957_/D __dut__._2661_/Y VGND VGND VPWR
+ VPWR __dut__._2957_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1908_ __dut__._2004_/A1 tie[106] __dut__._1907_/X VGND VGND VPWR VPWR __dut__._3011_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2888_ __dut__._3102_/CLK __dut__._2888_/D __dut__._2730_/Y VGND VGND VPWR
+ VPWR __dut__._2888_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1839_ __dut__._2507_/A __dut__._2976_/Q VGND VGND VPWR VPWR __dut__._1839_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_68_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2401__B prod[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1628__A2 mc[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_103_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1564__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1310_ __dut__.__uuf__._1309_/Y __dut__.__uuf__._1294_/X __dut__.__uuf__._1296_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1310_/X sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._2799__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2290_ __dut__.__uuf__._2291_/CLK __dut__._2360_/X __dut__.__uuf__._1276_/X
+ VGND VGND VPWR VPWR __dut__._2361_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_132_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1241_ __dut__._2377_/B __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1241_/X sky130_fd_sc_hd__or2_4
XFILLER_113_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1172_ __dut__.__uuf__._1175_/A VGND VGND VPWR VPWR __dut__.__uuf__._1172_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2811_ clkbuf_5_2_0_tck/X __dut__._2811_/D __dut__._2807_/Y VGND VGND VPWR
+ VPWR __dut__._2811_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1508_ __dut__.__uuf__._1550_/A VGND VGND VPWR VPWR __dut__.__uuf__._1508_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2742_ rst VGND VGND VPWR VPWR __dut__._2742_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1439_ __dut__.__uuf__._1457_/A VGND VGND VPWR VPWR __dut__.__uuf__._1439_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2673_ rst VGND VGND VPWR VPWR __dut__._2673_/Y sky130_fd_sc_hd__inv_2
X__dut__._1624_ __dut__._1374_/Y mc[7] __dut__._1623_/X VGND VGND VPWR VPWR __dut__._1624_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1555_ __dut__._2509_/A __dut__._2855_/Q VGND VGND VPWR VPWR __dut__._1555_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_89_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1486_ __dut__._1490_/A1 __dut__._1484_/X __dut__._1485_/X VGND VGND VPWR
+ VPWR __dut__._2837_/D sky130_fd_sc_hd__a21o_4
XFILLER_73_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2107_ __dut__._2407_/A __dut__._2107_/B VGND VGND VPWR VPWR __dut__._2107_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._3087_ __dut__._3109_/CLK __dut__._3087_/D __dut__._2531_/Y VGND VGND VPWR
+ VPWR __dut__._3087_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2038_ __dut__._2044_/A1 prod[1] __dut__._2037_/X VGND VGND VPWR VPWR __dut__._3076_/D
+ sky130_fd_sc_hd__a21o_4
X_296_ _315_/CLK _296_/D trst VGND VGND VPWR VPWR _296_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_13_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_220_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1790_ __dut__.__uuf__._1790_/A __dut__.__uuf__._1790_/B __dut__.__uuf__._1790_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1791_/A sky130_fd_sc_hd__or3_4
XFILLER_60_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2342_ __dut__.__uuf__._2353_/CLK __dut__._2464_/X __dut__.__uuf__._1093_/X
+ VGND VGND VPWR VPWR prod[41] sky130_fd_sc_hd__dfrtp_4
XFILLER_133_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2273_ __dut__.__uuf__._2278_/CLK __dut__._2326_/X __dut__.__uuf__._1367_/X
+ VGND VGND VPWR VPWR __dut__._2327_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_114_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1224_ __dut__._2379_/B __dut__.__uuf__._1240_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1227_/B sky130_fd_sc_hd__and2_4
XFILLER_87_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1155_ __dut__.__uuf__._1161_/A VGND VGND VPWR VPWR __dut__.__uuf__._1155_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1086_ __dut__.__uuf__._1072_/X __dut__.__uuf__._1085_/X prod[44]
+ prod[45] __dut__.__uuf__._1082_/X VGND VGND VPWR VPWR __dut__._2470_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._3010_ _274_/CLK __dut__._3010_/D __dut__._2608_/Y VGND VGND VPWR VPWR __dut__._3010_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1988_ __dut__._1616_/X __dut__.__uuf__._1988_/B VGND VGND VPWR VPWR
+ __dut__._2106_/A2 sky130_fd_sc_hd__and2_4
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_150_ _146_/Y _296_/Q _308_/Q _307_/Q _220_/A VGND VGND VPWR VPWR _307_/D sky130_fd_sc_hd__o32a_4
XANTENNA___dut__._1401__A __dut__._2189_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2843__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1528__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2993__CLK __dut__._3093_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2725_ rst VGND VGND VPWR VPWR __dut__._2725_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2656_ rst VGND VGND VPWR VPWR __dut__._2656_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1607_ __dut__._2509_/A __dut__._2868_/Q VGND VGND VPWR VPWR __dut__._1607_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_120_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2587_ rst VGND VGND VPWR VPWR __dut__._2587_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1538_ __dut__._1562_/A1 __dut__._1536_/X __dut__._1537_/X VGND VGND VPWR
+ VPWR __dut__._2850_/D sky130_fd_sc_hd__a21o_4
X__dut__._1469_ __dut__._2325_/A __dut__._2831_/Q VGND VGND VPWR VPWR __dut__._1469_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2407__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_279_ _194_/A _279_/D VGND VGND VPWR VPWR _279_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_268_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_170_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1981__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1911_ __dut__.__uuf__._1867_/X __dut__.__uuf__._1909_/B __dut__.__uuf__._1909_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1912_/C sky130_fd_sc_hd__o21a_4
XFILLER_37_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1842_ __dut__.__uuf__._1842_/A VGND VGND VPWR VPWR __dut__.__uuf__._1842_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2317__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1773_ __dut__.__uuf__._1773_/A VGND VGND VPWR VPWR __dut__._2156_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_138_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0___dut__.__uuf__.__clk_source__ clkbuf_2_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_133_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2325_ __dut__.__uuf__._2328_/CLK __dut__._2430_/X __dut__.__uuf__._1143_/X
+ VGND VGND VPWR VPWR prod[24] sky130_fd_sc_hd__dfrtp_4
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2510_ __dut__._1374_/Y clk __dut__._2509_/X VGND VGND VPWR VPWR __dut__._2510_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2256_ __dut__.__uuf__._2293_/CLK __dut__._2292_/X __dut__.__uuf__._1451_/X
+ VGND VGND VPWR VPWR __dut__._2293_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2187_ __dut__.__uuf__._2216_/CLK __dut__._2154_/X __dut__.__uuf__._1618_/X
+ VGND VGND VPWR VPWR __dut__._2155_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2441_ __dut__._2507_/A prod[29] VGND VGND VPWR VPWR __dut__._2441_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1207_ __dut__.__uuf__._1206_/X __dut__.__uuf__._1203_/X prod[3]
+ prod[4] __dut__.__uuf__._1200_/X VGND VGND VPWR VPWR __dut__._2388_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1138_ __dut__.__uuf__._1132_/X __dut__.__uuf__._1129_/X prod[26]
+ prod[27] __dut__.__uuf__._1126_/X VGND VGND VPWR VPWR __dut__._2434_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_68_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2372_ __dut__._2376_/A1 __dut__._2372_/A2 __dut__._2371_/X VGND VGND VPWR
+ VPWR __dut__._2372_/X sky130_fd_sc_hd__a21o_4
XFILLER_28_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1069_ __dut__.__uuf__._1099_/A VGND VGND VPWR VPWR __dut__.__uuf__._1069_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_28_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_202_ _203_/A VGND VGND VPWR VPWR _202_/X sky130_fd_sc_hd__buf_2
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2227__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3021__CLK clkbuf_opt_1_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_133_ _131_/Y _231_/A _132_/Y _128_/X VGND VGND VPWR VPWR _134_/A sky130_fd_sc_hd__a211o_4
XFILLER_137_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1033__B2 __dut__.__uuf__._1025_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2708_ rst VGND VGND VPWR VPWR __dut__._2708_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2639_ rst VGND VGND VPWR VPWR __dut__._2639_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2889__CLK __dut__._3102_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_20_0_tck clkbuf_5_21_0_tck/A VGND VGND VPWR VPWR __dut__._3102_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1695__B __dut__._2904_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1912__A1 __dut__._2004_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2110_ VGND VGND VPWR VPWR __dut__.__uuf__._2110_/HI tie[117] sky130_fd_sc_hd__conb_1
XFILLER_130_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2041_ VGND VGND VPWR VPWR __dut__.__uuf__._2041_/HI tie[48] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2600__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._3044__CLK __dut__._3058_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1825_ __dut__.__uuf__._1813_/X __dut__.__uuf__._1823_/B __dut__.__uuf__._1823_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1826_/C sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._2047__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1756_ __dut__._2151_/B __dut__._2157_/B __dut__.__uuf__._1755_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1757_/C sky130_fd_sc_hd__o21ai_4
XFILLER_138_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2990_ __dut__._3093_/CLK __dut__._2990_/D __dut__._2628_/Y VGND VGND VPWR
+ VPWR __dut__._2990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1687_ __dut__._1508_/X VGND VGND VPWR VPWR __dut__.__uuf__._1691_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._1941_ __dut__._2189_/A __dut__._3027_/Q VGND VGND VPWR VPWR __dut__._1941_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2156__A1 __dut__._2172_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1872_ __dut__._1872_/A1 tie[88] __dut__._1871_/X VGND VGND VPWR VPWR __dut__._2993_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2308_ __dut__.__uuf__._2334_/CLK __dut__._2396_/X __dut__.__uuf__._1195_/X
+ VGND VGND VPWR VPWR prod[7] sky130_fd_sc_hd__dfrtp_4
XFILLER_125_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2239_ __dut__.__uuf__._2240_/CLK __dut__._2258_/X __dut__.__uuf__._1522_/X
+ VGND VGND VPWR VPWR __dut__._2259_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2424_ __dut__._2424_/A1 __dut__._2424_/A2 __dut__._2423_/X VGND VGND VPWR
+ VPWR __dut__._2424_/X sky130_fd_sc_hd__a21o_4
XFILLER_141_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_71_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2355_ __dut__._2407_/A __dut__._2355_/B VGND VGND VPWR VPWR __dut__._2355_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2286_ __dut__._2288_/A1 __dut__._2286_/A2 __dut__._2285_/X VGND VGND VPWR
+ VPWR __dut__._2286_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1190__B1 prod[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3067__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_133_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2386__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2197__CLK __dut__.__uuf__._2230_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1610_ __dut__.__uuf__._1628_/A VGND VGND VPWR VPWR __dut__.__uuf__._1615_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_147_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1541_ __dut__._1500_/X __dut__.__uuf__._1529_/X __dut__._2253_/B
+ __dut__.__uuf__._1534_/X VGND VGND VPWR VPWR __dut__.__uuf__._1541_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1472_ __dut__.__uuf__._1463_/X __dut__.__uuf__._1458_/X __dut__._2285_/B
+ __dut__.__uuf__._1469_/X __dut__.__uuf__._1471_/X VGND VGND VPWR VPWR __dut__._2284_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_143_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2024_ VGND VGND VPWR VPWR __dut__.__uuf__._2024_/HI tie[31] sky130_fd_sc_hd__conb_1
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2140_ __dut__._2140_/A1 __dut__._2140_/A2 __dut__._2139_/X VGND VGND VPWR
+ VPWR __dut__._2140_/X sky130_fd_sc_hd__a21o_4
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2071_ __dut__._2071_/A __dut__._3092_/Q VGND VGND VPWR VPWR __dut__._2071_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__.__uuf__._1236__A1 __dut__.__uuf__._1214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1808_ __dut__._2171_/B __dut__._2177_/B VGND VGND VPWR VPWR __dut__.__uuf__._1809_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_139_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1739_ __dut__.__uuf__._1761_/A __dut__.__uuf__._1739_/B __dut__.__uuf__._1739_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1740_/A sky130_fd_sc_hd__or3_4
X__dut__._2973_ __dut__._2985_/CLK __dut__._2973_/D __dut__._2645_/Y VGND VGND VPWR
+ VPWR __dut__._2973_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1924_ __dut__._1924_/A1 tie[114] __dut__._1923_/X VGND VGND VPWR VPWR __dut__._3019_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1855_ __dut__._1881_/A __dut__._2984_/Q VGND VGND VPWR VPWR __dut__._1855_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1786_ __dut__._1786_/A1 tie[45] __dut__._1785_/X VGND VGND VPWR VPWR __dut__._2950_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_96_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_5_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2407_ __dut__._2407_/A prod[12] VGND VGND VPWR VPWR __dut__._2407_/X sky130_fd_sc_hd__and2_4
XFILLER_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2338_ __dut__._2368_/A1 __dut__._2338_/A2 __dut__._2337_/X VGND VGND VPWR
+ VPWR __dut__._2338_/X sky130_fd_sc_hd__a21o_4
XFILLER_45_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2269_ __dut__._2269_/A __dut__._2269_/B VGND VGND VPWR VPWR __dut__._2269_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xpsn_inst_psn_buff_220 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2429_/A sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2927__CLK clkbuf_5_9_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_231 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2037_/A sky130_fd_sc_hd__buf_2
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_242 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1787_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_264 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2263_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_253 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1609_/A sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2368__A1 __dut__._2368_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_286 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2281_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_275 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1437_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_297 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2503_/A sky130_fd_sc_hd__buf_2
XFILLER_129_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_250_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2325__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1524_ __dut__._1520_/X __dut__.__uuf__._1508_/X __dut__._2261_/B
+ __dut__.__uuf__._1513_/X VGND VGND VPWR VPWR __dut__.__uuf__._1524_/X sky130_fd_sc_hd__o22a_4
XFILLER_151_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1455_ __dut__._1588_/X __dut__.__uuf__._1442_/X __dut__._2293_/B
+ __dut__.__uuf__._1448_/X VGND VGND VPWR VPWR __dut__.__uuf__._1455_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__.__uuf__._1796__A __dut__.__uuf__._1904_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1386_ __dut__.__uuf__._1386_/A VGND VGND VPWR VPWR __dut__.__uuf__._1386_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1640_ __dut__._2502_/A1 prod[37] __dut__._1639_/X VGND VGND VPWR VPWR __dut__._2877_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2212__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_131_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1571_ __dut__._2509_/A __dut__._2859_/Q VGND VGND VPWR VPWR __dut__._1571_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_112_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2007_ VGND VGND VPWR VPWR __dut__.__uuf__._2007_/HI tie[14] sky130_fd_sc_hd__conb_1
XFILLER_122_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2123_ __dut__._2325_/A __dut__._2123_/B VGND VGND VPWR VPWR __dut__._2123_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1036__A __dut__.__uuf__._1214_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_34_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2054_ __dut__._2412_/A1 prod[9] __dut__._2053_/X VGND VGND VPWR VPWR __dut__._3084_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2235__A __dut__._2325_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2956_ __dut__._2985_/CLK __dut__._2956_/D __dut__._2662_/Y VGND VGND VPWR
+ VPWR __dut__._2956_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1907_ __dut__._2005_/A __dut__._3010_/Q VGND VGND VPWR VPWR __dut__._1907_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2887_ __dut__._3102_/CLK __dut__._2887_/D __dut__._2731_/Y VGND VGND VPWR
+ VPWR __dut__._2887_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1838_ __dut__._1838_/A1 tie[71] __dut__._1837_/X VGND VGND VPWR VPWR __dut__._2976_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_110_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1769_ __dut__._1775_/A __dut__._2941_/Q VGND VGND VPWR VPWR __dut__._1769_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3105__CLK __dut__._3106_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2145__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1564__A2 mp[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2235__CLK __dut__.__uuf__._2240_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_298_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_4_0___dut__.__uuf__.__clk_source__ clkbuf_4_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2216_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_99_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_13_0_tck clkbuf_3_6_0_tck/X VGND VGND VPWR VPWR clkbuf_5_27_0_tck/A sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1240_ __dut__.__uuf__._1240_/A VGND VGND VPWR VPWR __dut__.__uuf__._1240_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1171_ __dut__.__uuf__._1162_/X __dut__.__uuf__._1159_/X prod[15]
+ prod[16] __dut__.__uuf__._1170_/X VGND VGND VPWR VPWR __dut__._2412_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_113_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2055__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2810_ __dut__._2860_/CLK __dut__._2810_/D __dut__._2808_/Y VGND VGND VPWR
+ VPWR __dut__._2810_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1507_ __dut__.__uuf__._1549_/A VGND VGND VPWR VPWR __dut__.__uuf__._1507_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2741_ rst VGND VGND VPWR VPWR __dut__._2741_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2672_ rst VGND VGND VPWR VPWR __dut__._2672_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1438_ __dut__.__uuf__._1461_/A VGND VGND VPWR VPWR __dut__.__uuf__._1457_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1623_ __dut__._2509_/A __dut__._2872_/Q VGND VGND VPWR VPWR __dut__._1623_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1369_ __dut__.__uuf__._1368_/Y __dut__.__uuf__._1347_/X __dut__.__uuf__._1348_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1369_/X sky130_fd_sc_hd__o21a_4
XFILLER_133_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1127__B1 prod[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1554_ __dut__._1554_/A1 __dut__._1552_/X __dut__._1553_/X VGND VGND VPWR
+ VPWR __dut__._2854_/D sky130_fd_sc_hd__a21o_4
XFILLER_46_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1485_ __dut__._2281_/A __dut__._2836_/Q VGND VGND VPWR VPWR __dut__._1485_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_133_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2106_ __dut__._2376_/A1 __dut__._2106_/A2 __dut__._2105_/X VGND VGND VPWR
+ VPWR __dut__._2106_/X sky130_fd_sc_hd__a21o_4
X__dut__._3086_ __dut__._3109_/CLK __dut__._3086_/D __dut__._2532_/Y VGND VGND VPWR
+ VPWR __dut__._3086_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2037_ __dut__._2037_/A __dut__._3075_/Q VGND VGND VPWR VPWR __dut__._2037_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_295_ _315_/CLK _295_/D trst VGND VGND VPWR VPWR _295_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2939_ __dut__._2941_/CLK __dut__._2939_/D __dut__._2679_/Y VGND VGND VPWR
+ VPWR __dut__._2939_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_tck clkbuf_3_3_0_tck/A VGND VGND VPWR VPWR clkbuf_4_5_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1979__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_213_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2603__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2341_ __dut__.__uuf__._2358_/CLK __dut__._2462_/X __dut__.__uuf__._1095_/X
+ VGND VGND VPWR VPWR prod[40] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2272_ __dut__.__uuf__._2278_/CLK __dut__._2324_/X __dut__.__uuf__._1371_/X
+ VGND VGND VPWR VPWR __dut__._2325_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_99_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1223_ __dut__._2377_/B __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1240_/A sky130_fd_sc_hd__and2_4
XFILLER_87_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1154_ __dut__.__uuf__._1147_/X __dut__.__uuf__._1144_/X prod[21]
+ prod[22] __dut__.__uuf__._1141_/X VGND VGND VPWR VPWR __dut__._2424_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__.__uuf__._1109__B1 prod[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1085_ __dut__.__uuf__._1099_/A VGND VGND VPWR VPWR __dut__.__uuf__._1085_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1124__A3 prod[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__300__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1889__A __dut__._2491_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1987_ __dut__.__uuf__._1980_/A __dut__.__uuf__._1985_/B __dut__.__uuf__._1023_/X
+ VGND VGND VPWR VPWR __dut__._2234_/A2 sky130_fd_sc_hd__o21a_4
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1528__A2 mp[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2513__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2724_ rst VGND VGND VPWR VPWR __dut__._2724_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2655_ rst VGND VGND VPWR VPWR __dut__._2655_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2586_ rst VGND VGND VPWR VPWR __dut__._2586_/Y sky130_fd_sc_hd__inv_2
X__dut__._1606_ __dut__._1606_/A1 __dut__._1604_/X __dut__._1605_/X VGND VGND VPWR
+ VPWR __dut__._2867_/D sky130_fd_sc_hd__a21o_4
XFILLER_120_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1537_ __dut__._1557_/A __dut__._2849_/Q VGND VGND VPWR VPWR __dut__._1537_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1468_ __dut__._1374_/Y mc[30] __dut__._1467_/X VGND VGND VPWR VPWR __dut__._1468_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1464__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1399_ __dut__._2509_/A __dut__._2816_/Q VGND VGND VPWR VPWR __dut__._1399_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_27_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1799__A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._3069_ clkbuf_5_5_0_tck/X __dut__._3069_/D __dut__._2549_/Y VGND VGND VPWR
+ VPWR __dut__._3069_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2407__B prod[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_278_ _194_/A _278_/D VGND VGND VPWR VPWR _278_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_163_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1910_ __dut__.__uuf__._1910_/A VGND VGND VPWR VPWR __dut__.__uuf__._1912_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1841_ __dut__._2183_/B __dut__._2189_/B VGND VGND VPWR VPWR __dut__.__uuf__._1842_/A
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1772_ __dut__.__uuf__._1815_/A __dut__.__uuf__._1772_/B __dut__.__uuf__._1772_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1773_/A sky130_fd_sc_hd__or3_4
XFILLER_134_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2333__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2324_ __dut__.__uuf__._2328_/CLK __dut__._2428_/X __dut__.__uuf__._1146_/X
+ VGND VGND VPWR VPWR prod[23] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2255_ __dut__.__uuf__._2293_/CLK __dut__._2290_/X __dut__.__uuf__._1454_/X
+ VGND VGND VPWR VPWR __dut__._2291_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_114_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2186_ __dut__.__uuf__._2216_/CLK __dut__._2152_/X __dut__.__uuf__._1619_/X
+ VGND VGND VPWR VPWR __dut__._2153_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2440_ __dut__._2440_/A1 __dut__._2440_/A2 __dut__._2439_/X VGND VGND VPWR
+ VPWR __dut__._2440_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1206_ __dut__.__uuf__._1463_/A VGND VGND VPWR VPWR __dut__.__uuf__._1206_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_102_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1137_ __dut__.__uuf__._1146_/A VGND VGND VPWR VPWR __dut__.__uuf__._1137_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_114_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2371_ __dut__._2407_/A __dut__._2371_/B VGND VGND VPWR VPWR __dut__._2371_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1068_ __dut__.__uuf__._1071_/A VGND VGND VPWR VPWR __dut__.__uuf__._1068_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_83_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2810__CLK __dut__._2860_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_201_ _203_/A VGND VGND VPWR VPWR _201_/X sky130_fd_sc_hd__buf_2
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_132_ _313_/Q _231_/A VGND VGND VPWR VPWR _132_/Y sky130_fd_sc_hd__nor2_4
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__.__uuf__._1033__A2 __dut__.__uuf__._1023_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2707_ rst VGND VGND VPWR VPWR __dut__._2707_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__293__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2638_ rst VGND VGND VPWR VPWR __dut__._2638_/Y sky130_fd_sc_hd__inv_2
X__dut__._2569_ rst VGND VGND VPWR VPWR __dut__._2569_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2153__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_280_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2040_ VGND VGND VPWR VPWR __dut__.__uuf__._2040_/HI tie[47] sky130_fd_sc_hd__conb_1
XFILLER_111_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1676__A1 __dut__._2502_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2833__CLK __dut__._2860_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1428__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1824_ __dut__.__uuf__._1824_/A VGND VGND VPWR VPWR __dut__.__uuf__._1826_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1600__A1 __dut__._1374_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1755_ __dut__.__uuf__._1755_/A VGND VGND VPWR VPWR __dut__.__uuf__._1755_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1686_ __dut__.__uuf__._1921_/A VGND VGND VPWR VPWR __dut__.__uuf__._1736_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1940_ __dut__._1942_/A1 tie[122] __dut__._1939_/X VGND VGND VPWR VPWR __dut__._3027_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_146_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1871_ __dut__._1881_/A __dut__._2992_/Q VGND VGND VPWR VPWR __dut__._1871_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2063__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2307_ __dut__.__uuf__._2307_/CLK __dut__._2394_/X __dut__.__uuf__._1197_/X
+ VGND VGND VPWR VPWR prod[6] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2238_ __dut__.__uuf__._2240_/CLK __dut__._2256_/X __dut__.__uuf__._1527_/X
+ VGND VGND VPWR VPWR __dut__._2257_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_88_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2423_ __dut__._2423_/A prod[20] VGND VGND VPWR VPWR __dut__._2423_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1407__A __dut__._2509_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2169_ __dut__.__uuf__._2291_/CLK __dut__._2118_/X __dut__.__uuf__._1639_/X
+ VGND VGND VPWR VPWR __dut__._2119_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1039__A __dut__.__uuf__._1464_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2354_ __dut__._2368_/A1 __dut__._2354_/A2 __dut__._2353_/X VGND VGND VPWR
+ VPWR __dut__._2354_/X sky130_fd_sc_hd__a21o_4
XFILLER_141_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_64_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2285_ __dut__._2303_/A __dut__._2285_/B VGND VGND VPWR VPWR __dut__._2285_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1502__A __dut__.__uuf__._1563_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2701__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2856__CLK __dut__._2860_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1658__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_126_A __dut__._1418_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1987__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1540_ __dut__.__uuf__._1543_/A VGND VGND VPWR VPWR __dut__.__uuf__._1540_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1471_ __dut__._1576_/X __dut__.__uuf__._1465_/X __dut__._2287_/B
+ __dut__.__uuf__._1470_/X VGND VGND VPWR VPWR __dut__.__uuf__._1471_/X sky130_fd_sc_hd__o22a_4
XFILLER_155_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2611__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2023_ VGND VGND VPWR VPWR __dut__.__uuf__._2023_/HI tie[30] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._3011__CLK _274_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2070_ __dut__._2422_/A1 prod[17] __dut__._2069_/X VGND VGND VPWR VPWR __dut__._3092_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_80_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1897__A __dut__._2005_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1807_ __dut__._1396_/X VGND VGND VPWR VPWR __dut__.__uuf__._1811_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_40_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1738_ __dut__.__uuf__._1704_/X __dut__.__uuf__._1736_/B __dut__.__uuf__._1736_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1739_/C sky130_fd_sc_hd__o21a_4
X__dut__._2972_ __dut__._2985_/CLK __dut__._2972_/D __dut__._2646_/Y VGND VGND VPWR
+ VPWR __dut__._2972_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2505__B prod[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2291__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1923_ __dut__._2207_/A __dut__._3018_/Q VGND VGND VPWR VPWR __dut__._1923_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_107_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2879__CLK __dut__._3106_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1669_ __dut__._2119_/B __dut__._2125_/B __dut__.__uuf__._1668_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1670_/C sky130_fd_sc_hd__o21ai_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1888__A1 __dut__._2488_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1854_ __dut__._1864_/A1 tie[79] __dut__._1853_/X VGND VGND VPWR VPWR __dut__._2984_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2521__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1785_ __dut__._1785_/A __dut__._2949_/Q VGND VGND VPWR VPWR __dut__._1785_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1992__A __dut__.__uuf__._1992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2406_ __dut__._2412_/A1 __dut__._2406_/A2 __dut__._2405_/X VGND VGND VPWR
+ VPWR __dut__._2406_/X sky130_fd_sc_hd__a21o_4
XFILLER_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2337_ __dut__._2407_/A __dut__._2337_/B VGND VGND VPWR VPWR __dut__._2337_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2268_ __dut__._2268_/A1 __dut__._2268_/A2 __dut__._2267_/X VGND VGND VPWR
+ VPWR __dut__._2268_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_221 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2427_/A sky130_fd_sc_hd__buf_2
XFILLER_31_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_210 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2501_/A sky130_fd_sc_hd__buf_2
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_243 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1785_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_232 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2041_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_254 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2297_/A sky130_fd_sc_hd__buf_2
X__dut__._2199_ __dut__._2207_/A __dut__._2199_/B VGND VGND VPWR VPWR __dut__._2199_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_265 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._2261_/A sky130_fd_sc_hd__buf_2
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_287 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1565_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_276 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1441_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_298 __dut__._2507_/A VGND VGND VPWR VPWR __dut__._1891_/A sky130_fd_sc_hd__buf_2
XFILLER_129_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._3034__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_243_A __dut__._2507_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2164__CLK __dut__.__uuf__._2291_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2056__A1 __dut__._2412_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2606__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1523_ __dut__.__uuf__._1563_/A VGND VGND VPWR VPWR __dut__.__uuf__._1523_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1454_ __dut__.__uuf__._1457_/A VGND VGND VPWR VPWR __dut__.__uuf__._1454_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1385_ __dut__.__uuf__._1378_/X __dut__.__uuf__._1384_/X __dut__._2321_/B
+ __dut__.__uuf__._1378_/X VGND VGND VPWR VPWR __dut__._2320_/A2 sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._2341__A __dut__._2407_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1570_ __dut__._1570_/A1 __dut__._1568_/X __dut__._1569_/X VGND VGND VPWR
+ VPWR __dut__._2858_/D sky130_fd_sc_hd__a21o_4
XFILLER_106_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2006_ VGND VGND VPWR VPWR __dut__.__uuf__._2006_/HI tie[13] sky130_fd_sc_hd__conb_1
XFILLER_85_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2122_ __dut__._2332_/A1 __dut__._2122_/A2 __dut__._2121_/X VGND VGND VPWR
+ VPWR __dut__._2122_/X sky130_fd_sc_hd__a21o_4
XFILLER_81_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2053_ __dut__._2407_/A __dut__._3083_/Q VGND VGND VPWR VPWR __dut__._2053_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2516__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_27_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._3057__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2955_ __dut__._2958_/CLK __dut__._2955_/D __dut__._2663_/Y VGND VGND VPWR
+ VPWR __dut__._2955_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1906_ __dut__._2004_/A1 tie[105] __dut__._1905_/X VGND VGND VPWR VPWR __dut__._3010_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2886_ __dut__._3102_/CLK __dut__._2886_/D __dut__._2732_/Y VGND VGND VPWR
+ VPWR __dut__._2886_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1837_ __dut__._2507_/A __dut__._2975_/Q VGND VGND VPWR VPWR __dut__._1837_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_150_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2187__CLK __dut__.__uuf__._2216_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1768_ __dut__._1780_/A1 tie[36] __dut__._1767_/X VGND VGND VPWR VPWR __dut__._2941_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_102_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1699_ __dut__._2189_/A __dut__._2906_/Q VGND VGND VPWR VPWR __dut__._1699_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2161__A __dut__._2207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1170_ __dut__.__uuf__._1200_/A VGND VGND VPWR VPWR __dut__.__uuf__._1170_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_140_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

