magic
tech sky130A
magscale 1 2
timestamp 1612119374
<< obsli1 >>
rect 1104 2159 59219 57681
<< obsm1 >>
rect 1104 1300 59231 57712
<< metal2 >>
rect 15014 59200 15070 60000
rect 45006 59200 45062 60000
rect 7470 0 7526 800
rect 22466 0 22522 800
rect 37462 0 37518 800
rect 52458 0 52514 800
<< obsm2 >>
rect 3422 59144 14958 59673
rect 15126 59144 44950 59673
rect 45118 59144 59046 59673
rect 3422 856 59046 59144
rect 3422 167 7414 856
rect 7582 167 22410 856
rect 22578 167 37406 856
rect 37574 167 52402 856
rect 52570 167 59046 856
<< metal3 >>
rect 59200 59576 60000 59696
rect 59200 59168 60000 59288
rect 59200 58624 60000 58744
rect 59200 58216 60000 58336
rect 59200 57808 60000 57928
rect 59200 57264 60000 57384
rect 59200 56856 60000 56976
rect 59200 56448 60000 56568
rect 59200 55904 60000 56024
rect 59200 55496 60000 55616
rect 59200 54952 60000 55072
rect 59200 54544 60000 54664
rect 59200 54136 60000 54256
rect 59200 53592 60000 53712
rect 59200 53184 60000 53304
rect 59200 52776 60000 52896
rect 59200 52232 60000 52352
rect 59200 51824 60000 51944
rect 59200 51416 60000 51536
rect 59200 50872 60000 50992
rect 59200 50464 60000 50584
rect 59200 49920 60000 50040
rect 59200 49512 60000 49632
rect 59200 49104 60000 49224
rect 59200 48560 60000 48680
rect 59200 48152 60000 48272
rect 59200 47744 60000 47864
rect 59200 47200 60000 47320
rect 59200 46792 60000 46912
rect 59200 46384 60000 46504
rect 59200 45840 60000 45960
rect 59200 45432 60000 45552
rect 59200 44888 60000 45008
rect 59200 44480 60000 44600
rect 59200 44072 60000 44192
rect 59200 43528 60000 43648
rect 59200 43120 60000 43240
rect 59200 42712 60000 42832
rect 59200 42168 60000 42288
rect 59200 41760 60000 41880
rect 59200 41216 60000 41336
rect 59200 40808 60000 40928
rect 59200 40400 60000 40520
rect 59200 39856 60000 39976
rect 59200 39448 60000 39568
rect 59200 39040 60000 39160
rect 59200 38496 60000 38616
rect 59200 38088 60000 38208
rect 59200 37680 60000 37800
rect 59200 37136 60000 37256
rect 59200 36728 60000 36848
rect 59200 36184 60000 36304
rect 59200 35776 60000 35896
rect 59200 35368 60000 35488
rect 59200 34824 60000 34944
rect 59200 34416 60000 34536
rect 59200 34008 60000 34128
rect 59200 33464 60000 33584
rect 59200 33056 60000 33176
rect 59200 32648 60000 32768
rect 59200 32104 60000 32224
rect 59200 31696 60000 31816
rect 59200 31152 60000 31272
rect 59200 30744 60000 30864
rect 59200 30336 60000 30456
rect 0 29928 800 30048
rect 59200 29792 60000 29912
rect 59200 29384 60000 29504
rect 59200 28976 60000 29096
rect 59200 28432 60000 28552
rect 59200 28024 60000 28144
rect 59200 27480 60000 27600
rect 59200 27072 60000 27192
rect 59200 26664 60000 26784
rect 59200 26120 60000 26240
rect 59200 25712 60000 25832
rect 59200 25304 60000 25424
rect 59200 24760 60000 24880
rect 59200 24352 60000 24472
rect 59200 23944 60000 24064
rect 59200 23400 60000 23520
rect 59200 22992 60000 23112
rect 59200 22448 60000 22568
rect 59200 22040 60000 22160
rect 59200 21632 60000 21752
rect 59200 21088 60000 21208
rect 59200 20680 60000 20800
rect 59200 20272 60000 20392
rect 59200 19728 60000 19848
rect 59200 19320 60000 19440
rect 59200 18912 60000 19032
rect 59200 18368 60000 18488
rect 59200 17960 60000 18080
rect 59200 17416 60000 17536
rect 59200 17008 60000 17128
rect 59200 16600 60000 16720
rect 59200 16056 60000 16176
rect 59200 15648 60000 15768
rect 59200 15240 60000 15360
rect 59200 14696 60000 14816
rect 59200 14288 60000 14408
rect 59200 13744 60000 13864
rect 59200 13336 60000 13456
rect 59200 12928 60000 13048
rect 59200 12384 60000 12504
rect 59200 11976 60000 12096
rect 59200 11568 60000 11688
rect 59200 11024 60000 11144
rect 59200 10616 60000 10736
rect 59200 10208 60000 10328
rect 59200 9664 60000 9784
rect 59200 9256 60000 9376
rect 59200 8712 60000 8832
rect 59200 8304 60000 8424
rect 59200 7896 60000 8016
rect 59200 7352 60000 7472
rect 59200 6944 60000 7064
rect 59200 6536 60000 6656
rect 59200 5992 60000 6112
rect 59200 5584 60000 5704
rect 59200 5176 60000 5296
rect 59200 4632 60000 4752
rect 59200 4224 60000 4344
rect 59200 3680 60000 3800
rect 59200 3272 60000 3392
rect 59200 2864 60000 2984
rect 59200 2320 60000 2440
rect 59200 1912 60000 2032
rect 59200 1504 60000 1624
rect 59200 960 60000 1080
rect 59200 552 60000 672
rect 59200 144 60000 264
<< obsm3 >>
rect 800 59496 59120 59669
rect 800 59368 59200 59496
rect 800 59088 59120 59368
rect 800 58824 59200 59088
rect 800 58544 59120 58824
rect 800 58416 59200 58544
rect 800 58136 59120 58416
rect 800 58008 59200 58136
rect 800 57728 59120 58008
rect 800 57464 59200 57728
rect 800 57184 59120 57464
rect 800 57056 59200 57184
rect 800 56776 59120 57056
rect 800 56648 59200 56776
rect 800 56368 59120 56648
rect 800 56104 59200 56368
rect 800 55824 59120 56104
rect 800 55696 59200 55824
rect 800 55416 59120 55696
rect 800 55152 59200 55416
rect 800 54872 59120 55152
rect 800 54744 59200 54872
rect 800 54464 59120 54744
rect 800 54336 59200 54464
rect 800 54056 59120 54336
rect 800 53792 59200 54056
rect 800 53512 59120 53792
rect 800 53384 59200 53512
rect 800 53104 59120 53384
rect 800 52976 59200 53104
rect 800 52696 59120 52976
rect 800 52432 59200 52696
rect 800 52152 59120 52432
rect 800 52024 59200 52152
rect 800 51744 59120 52024
rect 800 51616 59200 51744
rect 800 51336 59120 51616
rect 800 51072 59200 51336
rect 800 50792 59120 51072
rect 800 50664 59200 50792
rect 800 50384 59120 50664
rect 800 50120 59200 50384
rect 800 49840 59120 50120
rect 800 49712 59200 49840
rect 800 49432 59120 49712
rect 800 49304 59200 49432
rect 800 49024 59120 49304
rect 800 48760 59200 49024
rect 800 48480 59120 48760
rect 800 48352 59200 48480
rect 800 48072 59120 48352
rect 800 47944 59200 48072
rect 800 47664 59120 47944
rect 800 47400 59200 47664
rect 800 47120 59120 47400
rect 800 46992 59200 47120
rect 800 46712 59120 46992
rect 800 46584 59200 46712
rect 800 46304 59120 46584
rect 800 46040 59200 46304
rect 800 45760 59120 46040
rect 800 45632 59200 45760
rect 800 45352 59120 45632
rect 800 45088 59200 45352
rect 800 44808 59120 45088
rect 800 44680 59200 44808
rect 800 44400 59120 44680
rect 800 44272 59200 44400
rect 800 43992 59120 44272
rect 800 43728 59200 43992
rect 800 43448 59120 43728
rect 800 43320 59200 43448
rect 800 43040 59120 43320
rect 800 42912 59200 43040
rect 800 42632 59120 42912
rect 800 42368 59200 42632
rect 800 42088 59120 42368
rect 800 41960 59200 42088
rect 800 41680 59120 41960
rect 800 41416 59200 41680
rect 800 41136 59120 41416
rect 800 41008 59200 41136
rect 800 40728 59120 41008
rect 800 40600 59200 40728
rect 800 40320 59120 40600
rect 800 40056 59200 40320
rect 800 39776 59120 40056
rect 800 39648 59200 39776
rect 800 39368 59120 39648
rect 800 39240 59200 39368
rect 800 38960 59120 39240
rect 800 38696 59200 38960
rect 800 38416 59120 38696
rect 800 38288 59200 38416
rect 800 38008 59120 38288
rect 800 37880 59200 38008
rect 800 37600 59120 37880
rect 800 37336 59200 37600
rect 800 37056 59120 37336
rect 800 36928 59200 37056
rect 800 36648 59120 36928
rect 800 36384 59200 36648
rect 800 36104 59120 36384
rect 800 35976 59200 36104
rect 800 35696 59120 35976
rect 800 35568 59200 35696
rect 800 35288 59120 35568
rect 800 35024 59200 35288
rect 800 34744 59120 35024
rect 800 34616 59200 34744
rect 800 34336 59120 34616
rect 800 34208 59200 34336
rect 800 33928 59120 34208
rect 800 33664 59200 33928
rect 800 33384 59120 33664
rect 800 33256 59200 33384
rect 800 32976 59120 33256
rect 800 32848 59200 32976
rect 800 32568 59120 32848
rect 800 32304 59200 32568
rect 800 32024 59120 32304
rect 800 31896 59200 32024
rect 800 31616 59120 31896
rect 800 31352 59200 31616
rect 800 31072 59120 31352
rect 800 30944 59200 31072
rect 800 30664 59120 30944
rect 800 30536 59200 30664
rect 800 30256 59120 30536
rect 800 30128 59200 30256
rect 880 29992 59200 30128
rect 880 29848 59120 29992
rect 800 29712 59120 29848
rect 800 29584 59200 29712
rect 800 29304 59120 29584
rect 800 29176 59200 29304
rect 800 28896 59120 29176
rect 800 28632 59200 28896
rect 800 28352 59120 28632
rect 800 28224 59200 28352
rect 800 27944 59120 28224
rect 800 27680 59200 27944
rect 800 27400 59120 27680
rect 800 27272 59200 27400
rect 800 26992 59120 27272
rect 800 26864 59200 26992
rect 800 26584 59120 26864
rect 800 26320 59200 26584
rect 800 26040 59120 26320
rect 800 25912 59200 26040
rect 800 25632 59120 25912
rect 800 25504 59200 25632
rect 800 25224 59120 25504
rect 800 24960 59200 25224
rect 800 24680 59120 24960
rect 800 24552 59200 24680
rect 800 24272 59120 24552
rect 800 24144 59200 24272
rect 800 23864 59120 24144
rect 800 23600 59200 23864
rect 800 23320 59120 23600
rect 800 23192 59200 23320
rect 800 22912 59120 23192
rect 800 22648 59200 22912
rect 800 22368 59120 22648
rect 800 22240 59200 22368
rect 800 21960 59120 22240
rect 800 21832 59200 21960
rect 800 21552 59120 21832
rect 800 21288 59200 21552
rect 800 21008 59120 21288
rect 800 20880 59200 21008
rect 800 20600 59120 20880
rect 800 20472 59200 20600
rect 800 20192 59120 20472
rect 800 19928 59200 20192
rect 800 19648 59120 19928
rect 800 19520 59200 19648
rect 800 19240 59120 19520
rect 800 19112 59200 19240
rect 800 18832 59120 19112
rect 800 18568 59200 18832
rect 800 18288 59120 18568
rect 800 18160 59200 18288
rect 800 17880 59120 18160
rect 800 17616 59200 17880
rect 800 17336 59120 17616
rect 800 17208 59200 17336
rect 800 16928 59120 17208
rect 800 16800 59200 16928
rect 800 16520 59120 16800
rect 800 16256 59200 16520
rect 800 15976 59120 16256
rect 800 15848 59200 15976
rect 800 15568 59120 15848
rect 800 15440 59200 15568
rect 800 15160 59120 15440
rect 800 14896 59200 15160
rect 800 14616 59120 14896
rect 800 14488 59200 14616
rect 800 14208 59120 14488
rect 800 13944 59200 14208
rect 800 13664 59120 13944
rect 800 13536 59200 13664
rect 800 13256 59120 13536
rect 800 13128 59200 13256
rect 800 12848 59120 13128
rect 800 12584 59200 12848
rect 800 12304 59120 12584
rect 800 12176 59200 12304
rect 800 11896 59120 12176
rect 800 11768 59200 11896
rect 800 11488 59120 11768
rect 800 11224 59200 11488
rect 800 10944 59120 11224
rect 800 10816 59200 10944
rect 800 10536 59120 10816
rect 800 10408 59200 10536
rect 800 10128 59120 10408
rect 800 9864 59200 10128
rect 800 9584 59120 9864
rect 800 9456 59200 9584
rect 800 9176 59120 9456
rect 800 8912 59200 9176
rect 800 8632 59120 8912
rect 800 8504 59200 8632
rect 800 8224 59120 8504
rect 800 8096 59200 8224
rect 800 7816 59120 8096
rect 800 7552 59200 7816
rect 800 7272 59120 7552
rect 800 7144 59200 7272
rect 800 6864 59120 7144
rect 800 6736 59200 6864
rect 800 6456 59120 6736
rect 800 6192 59200 6456
rect 800 5912 59120 6192
rect 800 5784 59200 5912
rect 800 5504 59120 5784
rect 800 5376 59200 5504
rect 800 5096 59120 5376
rect 800 4832 59200 5096
rect 800 4552 59120 4832
rect 800 4424 59200 4552
rect 800 4144 59120 4424
rect 800 3880 59200 4144
rect 800 3600 59120 3880
rect 800 3472 59200 3600
rect 800 3192 59120 3472
rect 800 3064 59200 3192
rect 800 2784 59120 3064
rect 800 2520 59200 2784
rect 800 2240 59120 2520
rect 800 2112 59200 2240
rect 800 1832 59120 2112
rect 800 1704 59200 1832
rect 800 1424 59120 1704
rect 800 1160 59200 1424
rect 800 880 59120 1160
rect 800 752 59200 880
rect 800 472 59120 752
rect 800 344 59200 472
rect 800 171 59120 344
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< labels >>
rlabel metal2 s 7470 0 7526 800 6 clk
port 1 nsew signal input
rlabel metal3 s 59200 59168 60000 59288 6 done
port 2 nsew signal output
rlabel metal3 s 59200 144 60000 264 6 mc[0]
port 3 nsew signal input
rlabel metal3 s 59200 4632 60000 4752 6 mc[10]
port 4 nsew signal input
rlabel metal3 s 59200 5176 60000 5296 6 mc[11]
port 5 nsew signal input
rlabel metal3 s 59200 5584 60000 5704 6 mc[12]
port 6 nsew signal input
rlabel metal3 s 59200 5992 60000 6112 6 mc[13]
port 7 nsew signal input
rlabel metal3 s 59200 6536 60000 6656 6 mc[14]
port 8 nsew signal input
rlabel metal3 s 59200 6944 60000 7064 6 mc[15]
port 9 nsew signal input
rlabel metal3 s 59200 7352 60000 7472 6 mc[16]
port 10 nsew signal input
rlabel metal3 s 59200 7896 60000 8016 6 mc[17]
port 11 nsew signal input
rlabel metal3 s 59200 8304 60000 8424 6 mc[18]
port 12 nsew signal input
rlabel metal3 s 59200 8712 60000 8832 6 mc[19]
port 13 nsew signal input
rlabel metal3 s 59200 552 60000 672 6 mc[1]
port 14 nsew signal input
rlabel metal3 s 59200 9256 60000 9376 6 mc[20]
port 15 nsew signal input
rlabel metal3 s 59200 9664 60000 9784 6 mc[21]
port 16 nsew signal input
rlabel metal3 s 59200 10208 60000 10328 6 mc[22]
port 17 nsew signal input
rlabel metal3 s 59200 10616 60000 10736 6 mc[23]
port 18 nsew signal input
rlabel metal3 s 59200 11024 60000 11144 6 mc[24]
port 19 nsew signal input
rlabel metal3 s 59200 11568 60000 11688 6 mc[25]
port 20 nsew signal input
rlabel metal3 s 59200 11976 60000 12096 6 mc[26]
port 21 nsew signal input
rlabel metal3 s 59200 12384 60000 12504 6 mc[27]
port 22 nsew signal input
rlabel metal3 s 59200 12928 60000 13048 6 mc[28]
port 23 nsew signal input
rlabel metal3 s 59200 13336 60000 13456 6 mc[29]
port 24 nsew signal input
rlabel metal3 s 59200 960 60000 1080 6 mc[2]
port 25 nsew signal input
rlabel metal3 s 59200 13744 60000 13864 6 mc[30]
port 26 nsew signal input
rlabel metal3 s 59200 14288 60000 14408 6 mc[31]
port 27 nsew signal input
rlabel metal3 s 59200 1504 60000 1624 6 mc[3]
port 28 nsew signal input
rlabel metal3 s 59200 1912 60000 2032 6 mc[4]
port 29 nsew signal input
rlabel metal3 s 59200 2320 60000 2440 6 mc[5]
port 30 nsew signal input
rlabel metal3 s 59200 2864 60000 2984 6 mc[6]
port 31 nsew signal input
rlabel metal3 s 59200 3272 60000 3392 6 mc[7]
port 32 nsew signal input
rlabel metal3 s 59200 3680 60000 3800 6 mc[8]
port 33 nsew signal input
rlabel metal3 s 59200 4224 60000 4344 6 mc[9]
port 34 nsew signal input
rlabel metal3 s 59200 14696 60000 14816 6 mp[0]
port 35 nsew signal input
rlabel metal3 s 59200 19320 60000 19440 6 mp[10]
port 36 nsew signal input
rlabel metal3 s 59200 19728 60000 19848 6 mp[11]
port 37 nsew signal input
rlabel metal3 s 59200 20272 60000 20392 6 mp[12]
port 38 nsew signal input
rlabel metal3 s 59200 20680 60000 20800 6 mp[13]
port 39 nsew signal input
rlabel metal3 s 59200 21088 60000 21208 6 mp[14]
port 40 nsew signal input
rlabel metal3 s 59200 21632 60000 21752 6 mp[15]
port 41 nsew signal input
rlabel metal3 s 59200 22040 60000 22160 6 mp[16]
port 42 nsew signal input
rlabel metal3 s 59200 22448 60000 22568 6 mp[17]
port 43 nsew signal input
rlabel metal3 s 59200 22992 60000 23112 6 mp[18]
port 44 nsew signal input
rlabel metal3 s 59200 23400 60000 23520 6 mp[19]
port 45 nsew signal input
rlabel metal3 s 59200 15240 60000 15360 6 mp[1]
port 46 nsew signal input
rlabel metal3 s 59200 23944 60000 24064 6 mp[20]
port 47 nsew signal input
rlabel metal3 s 59200 24352 60000 24472 6 mp[21]
port 48 nsew signal input
rlabel metal3 s 59200 24760 60000 24880 6 mp[22]
port 49 nsew signal input
rlabel metal3 s 59200 25304 60000 25424 6 mp[23]
port 50 nsew signal input
rlabel metal3 s 59200 25712 60000 25832 6 mp[24]
port 51 nsew signal input
rlabel metal3 s 59200 26120 60000 26240 6 mp[25]
port 52 nsew signal input
rlabel metal3 s 59200 26664 60000 26784 6 mp[26]
port 53 nsew signal input
rlabel metal3 s 59200 27072 60000 27192 6 mp[27]
port 54 nsew signal input
rlabel metal3 s 59200 27480 60000 27600 6 mp[28]
port 55 nsew signal input
rlabel metal3 s 59200 28024 60000 28144 6 mp[29]
port 56 nsew signal input
rlabel metal3 s 59200 15648 60000 15768 6 mp[2]
port 57 nsew signal input
rlabel metal3 s 59200 28432 60000 28552 6 mp[30]
port 58 nsew signal input
rlabel metal3 s 59200 28976 60000 29096 6 mp[31]
port 59 nsew signal input
rlabel metal3 s 59200 16056 60000 16176 6 mp[3]
port 60 nsew signal input
rlabel metal3 s 59200 16600 60000 16720 6 mp[4]
port 61 nsew signal input
rlabel metal3 s 59200 17008 60000 17128 6 mp[5]
port 62 nsew signal input
rlabel metal3 s 59200 17416 60000 17536 6 mp[6]
port 63 nsew signal input
rlabel metal3 s 59200 17960 60000 18080 6 mp[7]
port 64 nsew signal input
rlabel metal3 s 59200 18368 60000 18488 6 mp[8]
port 65 nsew signal input
rlabel metal3 s 59200 18912 60000 19032 6 mp[9]
port 66 nsew signal input
rlabel metal3 s 59200 29384 60000 29504 6 prod[0]
port 67 nsew signal output
rlabel metal3 s 59200 34008 60000 34128 6 prod[10]
port 68 nsew signal output
rlabel metal3 s 59200 34416 60000 34536 6 prod[11]
port 69 nsew signal output
rlabel metal3 s 59200 34824 60000 34944 6 prod[12]
port 70 nsew signal output
rlabel metal3 s 59200 35368 60000 35488 6 prod[13]
port 71 nsew signal output
rlabel metal3 s 59200 35776 60000 35896 6 prod[14]
port 72 nsew signal output
rlabel metal3 s 59200 36184 60000 36304 6 prod[15]
port 73 nsew signal output
rlabel metal3 s 59200 36728 60000 36848 6 prod[16]
port 74 nsew signal output
rlabel metal3 s 59200 37136 60000 37256 6 prod[17]
port 75 nsew signal output
rlabel metal3 s 59200 37680 60000 37800 6 prod[18]
port 76 nsew signal output
rlabel metal3 s 59200 38088 60000 38208 6 prod[19]
port 77 nsew signal output
rlabel metal3 s 59200 29792 60000 29912 6 prod[1]
port 78 nsew signal output
rlabel metal3 s 59200 38496 60000 38616 6 prod[20]
port 79 nsew signal output
rlabel metal3 s 59200 39040 60000 39160 6 prod[21]
port 80 nsew signal output
rlabel metal3 s 59200 39448 60000 39568 6 prod[22]
port 81 nsew signal output
rlabel metal3 s 59200 39856 60000 39976 6 prod[23]
port 82 nsew signal output
rlabel metal3 s 59200 40400 60000 40520 6 prod[24]
port 83 nsew signal output
rlabel metal3 s 59200 40808 60000 40928 6 prod[25]
port 84 nsew signal output
rlabel metal3 s 59200 41216 60000 41336 6 prod[26]
port 85 nsew signal output
rlabel metal3 s 59200 41760 60000 41880 6 prod[27]
port 86 nsew signal output
rlabel metal3 s 59200 42168 60000 42288 6 prod[28]
port 87 nsew signal output
rlabel metal3 s 59200 42712 60000 42832 6 prod[29]
port 88 nsew signal output
rlabel metal3 s 59200 30336 60000 30456 6 prod[2]
port 89 nsew signal output
rlabel metal3 s 59200 43120 60000 43240 6 prod[30]
port 90 nsew signal output
rlabel metal3 s 59200 43528 60000 43648 6 prod[31]
port 91 nsew signal output
rlabel metal3 s 59200 44072 60000 44192 6 prod[32]
port 92 nsew signal output
rlabel metal3 s 59200 44480 60000 44600 6 prod[33]
port 93 nsew signal output
rlabel metal3 s 59200 44888 60000 45008 6 prod[34]
port 94 nsew signal output
rlabel metal3 s 59200 45432 60000 45552 6 prod[35]
port 95 nsew signal output
rlabel metal3 s 59200 45840 60000 45960 6 prod[36]
port 96 nsew signal output
rlabel metal3 s 59200 46384 60000 46504 6 prod[37]
port 97 nsew signal output
rlabel metal3 s 59200 46792 60000 46912 6 prod[38]
port 98 nsew signal output
rlabel metal3 s 59200 47200 60000 47320 6 prod[39]
port 99 nsew signal output
rlabel metal3 s 59200 30744 60000 30864 6 prod[3]
port 100 nsew signal output
rlabel metal3 s 59200 47744 60000 47864 6 prod[40]
port 101 nsew signal output
rlabel metal3 s 59200 48152 60000 48272 6 prod[41]
port 102 nsew signal output
rlabel metal3 s 59200 48560 60000 48680 6 prod[42]
port 103 nsew signal output
rlabel metal3 s 59200 49104 60000 49224 6 prod[43]
port 104 nsew signal output
rlabel metal3 s 59200 49512 60000 49632 6 prod[44]
port 105 nsew signal output
rlabel metal3 s 59200 49920 60000 50040 6 prod[45]
port 106 nsew signal output
rlabel metal3 s 59200 50464 60000 50584 6 prod[46]
port 107 nsew signal output
rlabel metal3 s 59200 50872 60000 50992 6 prod[47]
port 108 nsew signal output
rlabel metal3 s 59200 51416 60000 51536 6 prod[48]
port 109 nsew signal output
rlabel metal3 s 59200 51824 60000 51944 6 prod[49]
port 110 nsew signal output
rlabel metal3 s 59200 31152 60000 31272 6 prod[4]
port 111 nsew signal output
rlabel metal3 s 59200 52232 60000 52352 6 prod[50]
port 112 nsew signal output
rlabel metal3 s 59200 52776 60000 52896 6 prod[51]
port 113 nsew signal output
rlabel metal3 s 59200 53184 60000 53304 6 prod[52]
port 114 nsew signal output
rlabel metal3 s 59200 53592 60000 53712 6 prod[53]
port 115 nsew signal output
rlabel metal3 s 59200 54136 60000 54256 6 prod[54]
port 116 nsew signal output
rlabel metal3 s 59200 54544 60000 54664 6 prod[55]
port 117 nsew signal output
rlabel metal3 s 59200 54952 60000 55072 6 prod[56]
port 118 nsew signal output
rlabel metal3 s 59200 55496 60000 55616 6 prod[57]
port 119 nsew signal output
rlabel metal3 s 59200 55904 60000 56024 6 prod[58]
port 120 nsew signal output
rlabel metal3 s 59200 56448 60000 56568 6 prod[59]
port 121 nsew signal output
rlabel metal3 s 59200 31696 60000 31816 6 prod[5]
port 122 nsew signal output
rlabel metal3 s 59200 56856 60000 56976 6 prod[60]
port 123 nsew signal output
rlabel metal3 s 59200 57264 60000 57384 6 prod[61]
port 124 nsew signal output
rlabel metal3 s 59200 57808 60000 57928 6 prod[62]
port 125 nsew signal output
rlabel metal3 s 59200 58216 60000 58336 6 prod[63]
port 126 nsew signal output
rlabel metal3 s 59200 32104 60000 32224 6 prod[6]
port 127 nsew signal output
rlabel metal3 s 59200 32648 60000 32768 6 prod[7]
port 128 nsew signal output
rlabel metal3 s 59200 33056 60000 33176 6 prod[8]
port 129 nsew signal output
rlabel metal3 s 59200 33464 60000 33584 6 prod[9]
port 130 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 rst
port 131 nsew signal input
rlabel metal3 s 59200 58624 60000 58744 6 start
port 132 nsew signal input
rlabel metal2 s 15014 59200 15070 60000 6 tck
port 133 nsew signal input
rlabel metal2 s 45006 59200 45062 60000 6 tdi
port 134 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 tdo
port 135 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 tdo_paden_o
port 136 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 tms
port 137 nsew signal input
rlabel metal3 s 59200 59576 60000 59696 6 trst
port 138 nsew signal input
rlabel metal4 s 34928 2128 35248 57712 6 VPWR
port 139 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 57712 6 VPWR
port 140 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 VGND
port 141 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 VGND
port 142 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60000 60000
string LEFview TRUE
string GDS_FILE /project/openlane/spm_top/runs/spm_top/results/magic/spm_top.gds
string GDS_END 7055716
string GDS_START 264176
<< end >>

