magic
tech sky130A
magscale 1 2
timestamp 1611915300
<< obsli1 >>
rect 1104 2159 59035 57681
<< obsm1 >>
rect 1104 1912 59050 57712
<< metal2 >>
rect 30010 59200 30066 60000
rect 5998 0 6054 800
rect 17958 0 18014 800
rect 29918 0 29974 800
rect 41970 0 42026 800
rect 53930 0 53986 800
<< obsm2 >>
rect 3054 59144 29954 59673
rect 30122 59144 59046 59673
rect 3054 856 59046 59144
rect 3054 167 5942 856
rect 6110 167 17902 856
rect 18070 167 29862 856
rect 30030 167 41914 856
rect 42082 167 53874 856
rect 54042 167 59046 856
<< metal3 >>
rect 59200 59576 60000 59696
rect 59200 59168 60000 59288
rect 59200 58624 60000 58744
rect 59200 58216 60000 58336
rect 59200 57808 60000 57928
rect 59200 57264 60000 57384
rect 59200 56856 60000 56976
rect 59200 56312 60000 56432
rect 59200 55904 60000 56024
rect 59200 55496 60000 55616
rect 59200 54952 60000 55072
rect 59200 54544 60000 54664
rect 59200 54000 60000 54120
rect 59200 53592 60000 53712
rect 59200 53184 60000 53304
rect 59200 52640 60000 52760
rect 59200 52232 60000 52352
rect 59200 51688 60000 51808
rect 59200 51280 60000 51400
rect 59200 50872 60000 50992
rect 59200 50328 60000 50448
rect 59200 49920 60000 50040
rect 59200 49376 60000 49496
rect 59200 48968 60000 49088
rect 59200 48560 60000 48680
rect 59200 48016 60000 48136
rect 59200 47608 60000 47728
rect 59200 47200 60000 47320
rect 59200 46656 60000 46776
rect 59200 46248 60000 46368
rect 59200 45704 60000 45824
rect 59200 45296 60000 45416
rect 0 44888 800 45008
rect 59200 44888 60000 45008
rect 59200 44344 60000 44464
rect 59200 43936 60000 44056
rect 59200 43392 60000 43512
rect 59200 42984 60000 43104
rect 59200 42576 60000 42696
rect 59200 42032 60000 42152
rect 59200 41624 60000 41744
rect 59200 41080 60000 41200
rect 59200 40672 60000 40792
rect 59200 40264 60000 40384
rect 59200 39720 60000 39840
rect 59200 39312 60000 39432
rect 59200 38768 60000 38888
rect 59200 38360 60000 38480
rect 59200 37952 60000 38072
rect 59200 37408 60000 37528
rect 59200 37000 60000 37120
rect 59200 36456 60000 36576
rect 59200 36048 60000 36168
rect 59200 35640 60000 35760
rect 59200 35096 60000 35216
rect 59200 34688 60000 34808
rect 59200 34280 60000 34400
rect 59200 33736 60000 33856
rect 59200 33328 60000 33448
rect 59200 32784 60000 32904
rect 59200 32376 60000 32496
rect 59200 31968 60000 32088
rect 59200 31424 60000 31544
rect 59200 31016 60000 31136
rect 59200 30472 60000 30592
rect 59200 30064 60000 30184
rect 59200 29656 60000 29776
rect 59200 29112 60000 29232
rect 59200 28704 60000 28824
rect 59200 28160 60000 28280
rect 59200 27752 60000 27872
rect 59200 27344 60000 27464
rect 59200 26800 60000 26920
rect 59200 26392 60000 26512
rect 59200 25848 60000 25968
rect 59200 25440 60000 25560
rect 59200 25032 60000 25152
rect 59200 24488 60000 24608
rect 59200 24080 60000 24200
rect 59200 23672 60000 23792
rect 59200 23128 60000 23248
rect 59200 22720 60000 22840
rect 59200 22176 60000 22296
rect 59200 21768 60000 21888
rect 59200 21360 60000 21480
rect 59200 20816 60000 20936
rect 59200 20408 60000 20528
rect 59200 19864 60000 19984
rect 59200 19456 60000 19576
rect 59200 19048 60000 19168
rect 59200 18504 60000 18624
rect 59200 18096 60000 18216
rect 59200 17552 60000 17672
rect 59200 17144 60000 17264
rect 59200 16736 60000 16856
rect 59200 16192 60000 16312
rect 59200 15784 60000 15904
rect 59200 15240 60000 15360
rect 0 14968 800 15088
rect 59200 14832 60000 14952
rect 59200 14424 60000 14544
rect 59200 13880 60000 14000
rect 59200 13472 60000 13592
rect 59200 12928 60000 13048
rect 59200 12520 60000 12640
rect 59200 12112 60000 12232
rect 59200 11568 60000 11688
rect 59200 11160 60000 11280
rect 59200 10752 60000 10872
rect 59200 10208 60000 10328
rect 59200 9800 60000 9920
rect 59200 9256 60000 9376
rect 59200 8848 60000 8968
rect 59200 8440 60000 8560
rect 59200 7896 60000 8016
rect 59200 7488 60000 7608
rect 59200 6944 60000 7064
rect 59200 6536 60000 6656
rect 59200 6128 60000 6248
rect 59200 5584 60000 5704
rect 59200 5176 60000 5296
rect 59200 4632 60000 4752
rect 59200 4224 60000 4344
rect 59200 3816 60000 3936
rect 59200 3272 60000 3392
rect 59200 2864 60000 2984
rect 59200 2320 60000 2440
rect 59200 1912 60000 2032
rect 59200 1504 60000 1624
rect 59200 960 60000 1080
rect 59200 552 60000 672
rect 59200 144 60000 264
<< obsm3 >>
rect 800 59496 59120 59669
rect 800 59368 59200 59496
rect 800 59088 59120 59368
rect 800 58824 59200 59088
rect 800 58544 59120 58824
rect 800 58416 59200 58544
rect 800 58136 59120 58416
rect 800 58008 59200 58136
rect 800 57728 59120 58008
rect 800 57464 59200 57728
rect 800 57184 59120 57464
rect 800 57056 59200 57184
rect 800 56776 59120 57056
rect 800 56512 59200 56776
rect 800 56232 59120 56512
rect 800 56104 59200 56232
rect 800 55824 59120 56104
rect 800 55696 59200 55824
rect 800 55416 59120 55696
rect 800 55152 59200 55416
rect 800 54872 59120 55152
rect 800 54744 59200 54872
rect 800 54464 59120 54744
rect 800 54200 59200 54464
rect 800 53920 59120 54200
rect 800 53792 59200 53920
rect 800 53512 59120 53792
rect 800 53384 59200 53512
rect 800 53104 59120 53384
rect 800 52840 59200 53104
rect 800 52560 59120 52840
rect 800 52432 59200 52560
rect 800 52152 59120 52432
rect 800 51888 59200 52152
rect 800 51608 59120 51888
rect 800 51480 59200 51608
rect 800 51200 59120 51480
rect 800 51072 59200 51200
rect 800 50792 59120 51072
rect 800 50528 59200 50792
rect 800 50248 59120 50528
rect 800 50120 59200 50248
rect 800 49840 59120 50120
rect 800 49576 59200 49840
rect 800 49296 59120 49576
rect 800 49168 59200 49296
rect 800 48888 59120 49168
rect 800 48760 59200 48888
rect 800 48480 59120 48760
rect 800 48216 59200 48480
rect 800 47936 59120 48216
rect 800 47808 59200 47936
rect 800 47528 59120 47808
rect 800 47400 59200 47528
rect 800 47120 59120 47400
rect 800 46856 59200 47120
rect 800 46576 59120 46856
rect 800 46448 59200 46576
rect 800 46168 59120 46448
rect 800 45904 59200 46168
rect 800 45624 59120 45904
rect 800 45496 59200 45624
rect 800 45216 59120 45496
rect 800 45088 59200 45216
rect 880 44808 59120 45088
rect 800 44544 59200 44808
rect 800 44264 59120 44544
rect 800 44136 59200 44264
rect 800 43856 59120 44136
rect 800 43592 59200 43856
rect 800 43312 59120 43592
rect 800 43184 59200 43312
rect 800 42904 59120 43184
rect 800 42776 59200 42904
rect 800 42496 59120 42776
rect 800 42232 59200 42496
rect 800 41952 59120 42232
rect 800 41824 59200 41952
rect 800 41544 59120 41824
rect 800 41280 59200 41544
rect 800 41000 59120 41280
rect 800 40872 59200 41000
rect 800 40592 59120 40872
rect 800 40464 59200 40592
rect 800 40184 59120 40464
rect 800 39920 59200 40184
rect 800 39640 59120 39920
rect 800 39512 59200 39640
rect 800 39232 59120 39512
rect 800 38968 59200 39232
rect 800 38688 59120 38968
rect 800 38560 59200 38688
rect 800 38280 59120 38560
rect 800 38152 59200 38280
rect 800 37872 59120 38152
rect 800 37608 59200 37872
rect 800 37328 59120 37608
rect 800 37200 59200 37328
rect 800 36920 59120 37200
rect 800 36656 59200 36920
rect 800 36376 59120 36656
rect 800 36248 59200 36376
rect 800 35968 59120 36248
rect 800 35840 59200 35968
rect 800 35560 59120 35840
rect 800 35296 59200 35560
rect 800 35016 59120 35296
rect 800 34888 59200 35016
rect 800 34608 59120 34888
rect 800 34480 59200 34608
rect 800 34200 59120 34480
rect 800 33936 59200 34200
rect 800 33656 59120 33936
rect 800 33528 59200 33656
rect 800 33248 59120 33528
rect 800 32984 59200 33248
rect 800 32704 59120 32984
rect 800 32576 59200 32704
rect 800 32296 59120 32576
rect 800 32168 59200 32296
rect 800 31888 59120 32168
rect 800 31624 59200 31888
rect 800 31344 59120 31624
rect 800 31216 59200 31344
rect 800 30936 59120 31216
rect 800 30672 59200 30936
rect 800 30392 59120 30672
rect 800 30264 59200 30392
rect 800 29984 59120 30264
rect 800 29856 59200 29984
rect 800 29576 59120 29856
rect 800 29312 59200 29576
rect 800 29032 59120 29312
rect 800 28904 59200 29032
rect 800 28624 59120 28904
rect 800 28360 59200 28624
rect 800 28080 59120 28360
rect 800 27952 59200 28080
rect 800 27672 59120 27952
rect 800 27544 59200 27672
rect 800 27264 59120 27544
rect 800 27000 59200 27264
rect 800 26720 59120 27000
rect 800 26592 59200 26720
rect 800 26312 59120 26592
rect 800 26048 59200 26312
rect 800 25768 59120 26048
rect 800 25640 59200 25768
rect 800 25360 59120 25640
rect 800 25232 59200 25360
rect 800 24952 59120 25232
rect 800 24688 59200 24952
rect 800 24408 59120 24688
rect 800 24280 59200 24408
rect 800 24000 59120 24280
rect 800 23872 59200 24000
rect 800 23592 59120 23872
rect 800 23328 59200 23592
rect 800 23048 59120 23328
rect 800 22920 59200 23048
rect 800 22640 59120 22920
rect 800 22376 59200 22640
rect 800 22096 59120 22376
rect 800 21968 59200 22096
rect 800 21688 59120 21968
rect 800 21560 59200 21688
rect 800 21280 59120 21560
rect 800 21016 59200 21280
rect 800 20736 59120 21016
rect 800 20608 59200 20736
rect 800 20328 59120 20608
rect 800 20064 59200 20328
rect 800 19784 59120 20064
rect 800 19656 59200 19784
rect 800 19376 59120 19656
rect 800 19248 59200 19376
rect 800 18968 59120 19248
rect 800 18704 59200 18968
rect 800 18424 59120 18704
rect 800 18296 59200 18424
rect 800 18016 59120 18296
rect 800 17752 59200 18016
rect 800 17472 59120 17752
rect 800 17344 59200 17472
rect 800 17064 59120 17344
rect 800 16936 59200 17064
rect 800 16656 59120 16936
rect 800 16392 59200 16656
rect 800 16112 59120 16392
rect 800 15984 59200 16112
rect 800 15704 59120 15984
rect 800 15440 59200 15704
rect 800 15168 59120 15440
rect 880 15160 59120 15168
rect 880 15032 59200 15160
rect 880 14888 59120 15032
rect 800 14752 59120 14888
rect 800 14624 59200 14752
rect 800 14344 59120 14624
rect 800 14080 59200 14344
rect 800 13800 59120 14080
rect 800 13672 59200 13800
rect 800 13392 59120 13672
rect 800 13128 59200 13392
rect 800 12848 59120 13128
rect 800 12720 59200 12848
rect 800 12440 59120 12720
rect 800 12312 59200 12440
rect 800 12032 59120 12312
rect 800 11768 59200 12032
rect 800 11488 59120 11768
rect 800 11360 59200 11488
rect 800 11080 59120 11360
rect 800 10952 59200 11080
rect 800 10672 59120 10952
rect 800 10408 59200 10672
rect 800 10128 59120 10408
rect 800 10000 59200 10128
rect 800 9720 59120 10000
rect 800 9456 59200 9720
rect 800 9176 59120 9456
rect 800 9048 59200 9176
rect 800 8768 59120 9048
rect 800 8640 59200 8768
rect 800 8360 59120 8640
rect 800 8096 59200 8360
rect 800 7816 59120 8096
rect 800 7688 59200 7816
rect 800 7408 59120 7688
rect 800 7144 59200 7408
rect 800 6864 59120 7144
rect 800 6736 59200 6864
rect 800 6456 59120 6736
rect 800 6328 59200 6456
rect 800 6048 59120 6328
rect 800 5784 59200 6048
rect 800 5504 59120 5784
rect 800 5376 59200 5504
rect 800 5096 59120 5376
rect 800 4832 59200 5096
rect 800 4552 59120 4832
rect 800 4424 59200 4552
rect 800 4144 59120 4424
rect 800 4016 59200 4144
rect 800 3736 59120 4016
rect 800 3472 59200 3736
rect 800 3192 59120 3472
rect 800 3064 59200 3192
rect 800 2784 59120 3064
rect 800 2520 59200 2784
rect 800 2240 59120 2520
rect 800 2112 59200 2240
rect 800 1832 59120 2112
rect 800 1704 59200 1832
rect 800 1424 59120 1704
rect 800 1160 59200 1424
rect 800 880 59120 1160
rect 800 752 59200 880
rect 800 472 59120 752
rect 800 344 59200 472
rect 800 171 59120 344
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< obsm4 >>
rect 55811 53891 55877 54773
<< labels >>
rlabel metal2 s 5998 0 6054 800 6 clk
port 1 nsew signal input
rlabel metal3 s 59200 59576 60000 59696 6 done
port 2 nsew signal output
rlabel metal3 s 59200 144 60000 264 6 mc[0]
port 3 nsew signal input
rlabel metal3 s 59200 4632 60000 4752 6 mc[10]
port 4 nsew signal input
rlabel metal3 s 59200 5176 60000 5296 6 mc[11]
port 5 nsew signal input
rlabel metal3 s 59200 5584 60000 5704 6 mc[12]
port 6 nsew signal input
rlabel metal3 s 59200 6128 60000 6248 6 mc[13]
port 7 nsew signal input
rlabel metal3 s 59200 6536 60000 6656 6 mc[14]
port 8 nsew signal input
rlabel metal3 s 59200 6944 60000 7064 6 mc[15]
port 9 nsew signal input
rlabel metal3 s 59200 7488 60000 7608 6 mc[16]
port 10 nsew signal input
rlabel metal3 s 59200 7896 60000 8016 6 mc[17]
port 11 nsew signal input
rlabel metal3 s 59200 8440 60000 8560 6 mc[18]
port 12 nsew signal input
rlabel metal3 s 59200 8848 60000 8968 6 mc[19]
port 13 nsew signal input
rlabel metal3 s 59200 552 60000 672 6 mc[1]
port 14 nsew signal input
rlabel metal3 s 59200 9256 60000 9376 6 mc[20]
port 15 nsew signal input
rlabel metal3 s 59200 9800 60000 9920 6 mc[21]
port 16 nsew signal input
rlabel metal3 s 59200 10208 60000 10328 6 mc[22]
port 17 nsew signal input
rlabel metal3 s 59200 10752 60000 10872 6 mc[23]
port 18 nsew signal input
rlabel metal3 s 59200 11160 60000 11280 6 mc[24]
port 19 nsew signal input
rlabel metal3 s 59200 11568 60000 11688 6 mc[25]
port 20 nsew signal input
rlabel metal3 s 59200 12112 60000 12232 6 mc[26]
port 21 nsew signal input
rlabel metal3 s 59200 12520 60000 12640 6 mc[27]
port 22 nsew signal input
rlabel metal3 s 59200 12928 60000 13048 6 mc[28]
port 23 nsew signal input
rlabel metal3 s 59200 13472 60000 13592 6 mc[29]
port 24 nsew signal input
rlabel metal3 s 59200 960 60000 1080 6 mc[2]
port 25 nsew signal input
rlabel metal3 s 59200 13880 60000 14000 6 mc[30]
port 26 nsew signal input
rlabel metal3 s 59200 14424 60000 14544 6 mc[31]
port 27 nsew signal input
rlabel metal3 s 59200 1504 60000 1624 6 mc[3]
port 28 nsew signal input
rlabel metal3 s 59200 1912 60000 2032 6 mc[4]
port 29 nsew signal input
rlabel metal3 s 59200 2320 60000 2440 6 mc[5]
port 30 nsew signal input
rlabel metal3 s 59200 2864 60000 2984 6 mc[6]
port 31 nsew signal input
rlabel metal3 s 59200 3272 60000 3392 6 mc[7]
port 32 nsew signal input
rlabel metal3 s 59200 3816 60000 3936 6 mc[8]
port 33 nsew signal input
rlabel metal3 s 59200 4224 60000 4344 6 mc[9]
port 34 nsew signal input
rlabel metal3 s 59200 14832 60000 14952 6 mp[0]
port 35 nsew signal input
rlabel metal3 s 59200 19456 60000 19576 6 mp[10]
port 36 nsew signal input
rlabel metal3 s 59200 19864 60000 19984 6 mp[11]
port 37 nsew signal input
rlabel metal3 s 59200 20408 60000 20528 6 mp[12]
port 38 nsew signal input
rlabel metal3 s 59200 20816 60000 20936 6 mp[13]
port 39 nsew signal input
rlabel metal3 s 59200 21360 60000 21480 6 mp[14]
port 40 nsew signal input
rlabel metal3 s 59200 21768 60000 21888 6 mp[15]
port 41 nsew signal input
rlabel metal3 s 59200 22176 60000 22296 6 mp[16]
port 42 nsew signal input
rlabel metal3 s 59200 22720 60000 22840 6 mp[17]
port 43 nsew signal input
rlabel metal3 s 59200 23128 60000 23248 6 mp[18]
port 44 nsew signal input
rlabel metal3 s 59200 23672 60000 23792 6 mp[19]
port 45 nsew signal input
rlabel metal3 s 59200 15240 60000 15360 6 mp[1]
port 46 nsew signal input
rlabel metal3 s 59200 24080 60000 24200 6 mp[20]
port 47 nsew signal input
rlabel metal3 s 59200 24488 60000 24608 6 mp[21]
port 48 nsew signal input
rlabel metal3 s 59200 25032 60000 25152 6 mp[22]
port 49 nsew signal input
rlabel metal3 s 59200 25440 60000 25560 6 mp[23]
port 50 nsew signal input
rlabel metal3 s 59200 25848 60000 25968 6 mp[24]
port 51 nsew signal input
rlabel metal3 s 59200 26392 60000 26512 6 mp[25]
port 52 nsew signal input
rlabel metal3 s 59200 26800 60000 26920 6 mp[26]
port 53 nsew signal input
rlabel metal3 s 59200 27344 60000 27464 6 mp[27]
port 54 nsew signal input
rlabel metal3 s 59200 27752 60000 27872 6 mp[28]
port 55 nsew signal input
rlabel metal3 s 59200 28160 60000 28280 6 mp[29]
port 56 nsew signal input
rlabel metal3 s 59200 15784 60000 15904 6 mp[2]
port 57 nsew signal input
rlabel metal3 s 59200 28704 60000 28824 6 mp[30]
port 58 nsew signal input
rlabel metal3 s 59200 29112 60000 29232 6 mp[31]
port 59 nsew signal input
rlabel metal3 s 59200 16192 60000 16312 6 mp[3]
port 60 nsew signal input
rlabel metal3 s 59200 16736 60000 16856 6 mp[4]
port 61 nsew signal input
rlabel metal3 s 59200 17144 60000 17264 6 mp[5]
port 62 nsew signal input
rlabel metal3 s 59200 17552 60000 17672 6 mp[6]
port 63 nsew signal input
rlabel metal3 s 59200 18096 60000 18216 6 mp[7]
port 64 nsew signal input
rlabel metal3 s 59200 18504 60000 18624 6 mp[8]
port 65 nsew signal input
rlabel metal3 s 59200 19048 60000 19168 6 mp[9]
port 66 nsew signal input
rlabel metal3 s 59200 29656 60000 29776 6 prod[0]
port 67 nsew signal output
rlabel metal3 s 59200 34280 60000 34400 6 prod[10]
port 68 nsew signal output
rlabel metal3 s 59200 34688 60000 34808 6 prod[11]
port 69 nsew signal output
rlabel metal3 s 59200 35096 60000 35216 6 prod[12]
port 70 nsew signal output
rlabel metal3 s 59200 35640 60000 35760 6 prod[13]
port 71 nsew signal output
rlabel metal3 s 59200 36048 60000 36168 6 prod[14]
port 72 nsew signal output
rlabel metal3 s 59200 36456 60000 36576 6 prod[15]
port 73 nsew signal output
rlabel metal3 s 59200 37000 60000 37120 6 prod[16]
port 74 nsew signal output
rlabel metal3 s 59200 37408 60000 37528 6 prod[17]
port 75 nsew signal output
rlabel metal3 s 59200 37952 60000 38072 6 prod[18]
port 76 nsew signal output
rlabel metal3 s 59200 38360 60000 38480 6 prod[19]
port 77 nsew signal output
rlabel metal3 s 59200 30064 60000 30184 6 prod[1]
port 78 nsew signal output
rlabel metal3 s 59200 38768 60000 38888 6 prod[20]
port 79 nsew signal output
rlabel metal3 s 59200 39312 60000 39432 6 prod[21]
port 80 nsew signal output
rlabel metal3 s 59200 39720 60000 39840 6 prod[22]
port 81 nsew signal output
rlabel metal3 s 59200 40264 60000 40384 6 prod[23]
port 82 nsew signal output
rlabel metal3 s 59200 40672 60000 40792 6 prod[24]
port 83 nsew signal output
rlabel metal3 s 59200 41080 60000 41200 6 prod[25]
port 84 nsew signal output
rlabel metal3 s 59200 41624 60000 41744 6 prod[26]
port 85 nsew signal output
rlabel metal3 s 59200 42032 60000 42152 6 prod[27]
port 86 nsew signal output
rlabel metal3 s 59200 42576 60000 42696 6 prod[28]
port 87 nsew signal output
rlabel metal3 s 59200 42984 60000 43104 6 prod[29]
port 88 nsew signal output
rlabel metal3 s 59200 30472 60000 30592 6 prod[2]
port 89 nsew signal output
rlabel metal3 s 59200 43392 60000 43512 6 prod[30]
port 90 nsew signal output
rlabel metal3 s 59200 43936 60000 44056 6 prod[31]
port 91 nsew signal output
rlabel metal3 s 59200 44344 60000 44464 6 prod[32]
port 92 nsew signal output
rlabel metal3 s 59200 44888 60000 45008 6 prod[33]
port 93 nsew signal output
rlabel metal3 s 59200 45296 60000 45416 6 prod[34]
port 94 nsew signal output
rlabel metal3 s 59200 45704 60000 45824 6 prod[35]
port 95 nsew signal output
rlabel metal3 s 59200 46248 60000 46368 6 prod[36]
port 96 nsew signal output
rlabel metal3 s 59200 46656 60000 46776 6 prod[37]
port 97 nsew signal output
rlabel metal3 s 59200 47200 60000 47320 6 prod[38]
port 98 nsew signal output
rlabel metal3 s 59200 47608 60000 47728 6 prod[39]
port 99 nsew signal output
rlabel metal3 s 59200 31016 60000 31136 6 prod[3]
port 100 nsew signal output
rlabel metal3 s 59200 48016 60000 48136 6 prod[40]
port 101 nsew signal output
rlabel metal3 s 59200 48560 60000 48680 6 prod[41]
port 102 nsew signal output
rlabel metal3 s 59200 48968 60000 49088 6 prod[42]
port 103 nsew signal output
rlabel metal3 s 59200 49376 60000 49496 6 prod[43]
port 104 nsew signal output
rlabel metal3 s 59200 49920 60000 50040 6 prod[44]
port 105 nsew signal output
rlabel metal3 s 59200 50328 60000 50448 6 prod[45]
port 106 nsew signal output
rlabel metal3 s 59200 50872 60000 50992 6 prod[46]
port 107 nsew signal output
rlabel metal3 s 59200 51280 60000 51400 6 prod[47]
port 108 nsew signal output
rlabel metal3 s 59200 51688 60000 51808 6 prod[48]
port 109 nsew signal output
rlabel metal3 s 59200 52232 60000 52352 6 prod[49]
port 110 nsew signal output
rlabel metal3 s 59200 31424 60000 31544 6 prod[4]
port 111 nsew signal output
rlabel metal3 s 59200 52640 60000 52760 6 prod[50]
port 112 nsew signal output
rlabel metal3 s 59200 53184 60000 53304 6 prod[51]
port 113 nsew signal output
rlabel metal3 s 59200 53592 60000 53712 6 prod[52]
port 114 nsew signal output
rlabel metal3 s 59200 54000 60000 54120 6 prod[53]
port 115 nsew signal output
rlabel metal3 s 59200 54544 60000 54664 6 prod[54]
port 116 nsew signal output
rlabel metal3 s 59200 54952 60000 55072 6 prod[55]
port 117 nsew signal output
rlabel metal3 s 59200 55496 60000 55616 6 prod[56]
port 118 nsew signal output
rlabel metal3 s 59200 55904 60000 56024 6 prod[57]
port 119 nsew signal output
rlabel metal3 s 59200 56312 60000 56432 6 prod[58]
port 120 nsew signal output
rlabel metal3 s 59200 56856 60000 56976 6 prod[59]
port 121 nsew signal output
rlabel metal3 s 59200 31968 60000 32088 6 prod[5]
port 122 nsew signal output
rlabel metal3 s 59200 57264 60000 57384 6 prod[60]
port 123 nsew signal output
rlabel metal3 s 59200 57808 60000 57928 6 prod[61]
port 124 nsew signal output
rlabel metal3 s 59200 58216 60000 58336 6 prod[62]
port 125 nsew signal output
rlabel metal3 s 59200 58624 60000 58744 6 prod[63]
port 126 nsew signal output
rlabel metal3 s 59200 32376 60000 32496 6 prod[6]
port 127 nsew signal output
rlabel metal3 s 59200 32784 60000 32904 6 prod[7]
port 128 nsew signal output
rlabel metal3 s 59200 33328 60000 33448 6 prod[8]
port 129 nsew signal output
rlabel metal3 s 59200 33736 60000 33856 6 prod[9]
port 130 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 rst
port 131 nsew signal input
rlabel metal3 s 59200 59168 60000 59288 6 start
port 132 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 tck
port 133 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 tdi
port 134 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 tdo
port 135 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 tdo_paden_o
port 136 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 tms
port 137 nsew signal input
rlabel metal2 s 30010 59200 30066 60000 6 trst
port 138 nsew signal input
rlabel metal4 s 34928 2128 35248 57712 6 VPWR
port 139 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 57712 6 VPWR
port 140 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 VGND
port 141 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 VGND
port 142 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60000 60000
string LEFview TRUE
string GDS_FILE /project/openlane/spm_top/runs/spm_top/results/magic/spm_top.gds
string GDS_END 6551218
string GDS_START 264176
<< end >>

