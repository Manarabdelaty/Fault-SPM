magic
tech sky130A
magscale 1 2
timestamp 1612364373
<< locali >>
rect 249073 327947 249107 328049
rect 279433 327811 279467 328117
rect 315865 327879 315899 328049
rect 317521 327607 317555 327913
rect 248613 323663 248647 325873
rect 127633 3383 127667 4097
rect 248889 3723 248923 3961
rect 311173 3927 311207 4097
rect 311265 3723 311299 3893
rect 248981 3587 249015 3689
rect 311357 3587 311391 3689
rect 311449 3315 311483 3553
<< viali >>
rect 279433 328117 279467 328151
rect 249073 328049 249107 328083
rect 249073 327913 249107 327947
rect 315865 328049 315899 328083
rect 315865 327845 315899 327879
rect 317521 327913 317555 327947
rect 279433 327777 279467 327811
rect 317521 327573 317555 327607
rect 248613 325873 248647 325907
rect 248613 323629 248647 323663
rect 127633 4097 127667 4131
rect 311173 4097 311207 4131
rect 248889 3961 248923 3995
rect 311173 3893 311207 3927
rect 311265 3893 311299 3927
rect 248889 3689 248923 3723
rect 248981 3689 249015 3723
rect 311265 3689 311299 3723
rect 311357 3689 311391 3723
rect 248981 3553 249015 3587
rect 311357 3553 311391 3587
rect 311449 3553 311483 3587
rect 127633 3349 127667 3383
rect 311449 3281 311483 3315
<< metal1 >>
rect 256602 700408 256608 700460
rect 256660 700448 256666 700460
rect 348786 700448 348792 700460
rect 256660 700420 348792 700448
rect 256660 700408 256666 700420
rect 348786 700408 348792 700420
rect 348844 700408 348850 700460
rect 251082 700340 251088 700392
rect 251140 700380 251146 700392
rect 413646 700380 413652 700392
rect 251140 700352 413652 700380
rect 251140 700340 251146 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 291102 700272 291108 700324
rect 291160 700312 291166 700324
rect 462314 700312 462320 700324
rect 291160 700284 462320 700312
rect 291160 700272 291166 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 331214 697552 331220 697604
rect 331272 697592 331278 697604
rect 332502 697592 332508 697604
rect 331272 697564 332508 697592
rect 331272 697552 331278 697564
rect 332502 697552 332508 697564
rect 332560 697552 332566 697604
rect 284938 696940 284944 696992
rect 284996 696980 285002 696992
rect 580166 696980 580172 696992
rect 284996 696952 580172 696980
rect 284996 696940 285002 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 14458 667944 14464 667956
rect 3476 667916 14464 667944
rect 3476 667904 3482 667916
rect 14458 667904 14464 667916
rect 14516 667904 14522 667956
rect 338758 650020 338764 650072
rect 338816 650060 338822 650072
rect 580166 650060 580172 650072
rect 338816 650032 580172 650060
rect 338816 650020 338822 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 393958 603100 393964 603152
rect 394016 603140 394022 603152
rect 580166 603140 580172 603152
rect 394016 603112 580172 603140
rect 394016 603100 394022 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 384298 556180 384304 556232
rect 384356 556220 384362 556232
rect 579798 556220 579804 556232
rect 384356 556192 579804 556220
rect 384356 556180 384362 556192
rect 579798 556180 579804 556192
rect 579856 556180 579862 556232
rect 3326 552032 3332 552084
rect 3384 552072 3390 552084
rect 19978 552072 19984 552084
rect 3384 552044 19984 552072
rect 3384 552032 3390 552044
rect 19978 552032 19984 552044
rect 20036 552032 20042 552084
rect 391198 545096 391204 545148
rect 391256 545136 391262 545148
rect 580166 545136 580172 545148
rect 391256 545108 580172 545136
rect 391256 545096 391262 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 380158 509260 380164 509312
rect 380216 509300 380222 509312
rect 579798 509300 579804 509312
rect 380216 509272 579804 509300
rect 380216 509260 380222 509272
rect 579798 509260 579804 509272
rect 579856 509260 579862 509312
rect 388438 498176 388444 498228
rect 388496 498216 388502 498228
rect 580166 498216 580172 498228
rect 388496 498188 580172 498216
rect 388496 498176 388502 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 395338 462340 395344 462392
rect 395396 462380 395402 462392
rect 579798 462380 579804 462392
rect 395396 462352 579804 462380
rect 395396 462340 395402 462352
rect 579798 462340 579804 462352
rect 579856 462340 579862 462392
rect 3142 437452 3148 437504
rect 3200 437492 3206 437504
rect 21358 437492 21364 437504
rect 3200 437464 21364 437492
rect 3200 437452 3206 437464
rect 21358 437452 21364 437464
rect 21416 437452 21422 437504
rect 282270 424940 282276 424992
rect 282328 424980 282334 424992
rect 284938 424980 284944 424992
rect 282328 424952 284944 424980
rect 282328 424940 282334 424952
rect 284938 424940 284944 424952
rect 284996 424940 285002 424992
rect 3142 423648 3148 423700
rect 3200 423688 3206 423700
rect 6178 423688 6184 423700
rect 3200 423660 6184 423688
rect 3200 423648 3206 423660
rect 6178 423648 6184 423660
rect 6236 423648 6242 423700
rect 260006 423512 260012 423564
rect 260064 423552 260070 423564
rect 282914 423552 282920 423564
rect 260064 423524 282920 423552
rect 260064 423512 260070 423524
rect 282914 423512 282920 423524
rect 282972 423512 282978 423564
rect 219342 423444 219348 423496
rect 219400 423484 219406 423496
rect 264422 423484 264428 423496
rect 219400 423456 264428 423484
rect 219400 423444 219406 423456
rect 264422 423444 264428 423456
rect 264480 423444 264486 423496
rect 267642 423444 267648 423496
rect 267700 423484 267706 423496
rect 304442 423484 304448 423496
rect 267700 423456 304448 423484
rect 267700 423444 267706 423456
rect 304442 423444 304448 423456
rect 304500 423444 304506 423496
rect 202782 423376 202788 423428
rect 202840 423416 202846 423428
rect 308950 423416 308956 423428
rect 202840 423388 308956 423416
rect 202840 423376 202846 423388
rect 308950 423376 308956 423388
rect 309008 423376 309014 423428
rect 154482 423308 154488 423360
rect 154540 423348 154546 423360
rect 268930 423348 268936 423360
rect 154540 423320 268936 423348
rect 154540 423308 154546 423320
rect 268930 423308 268936 423320
rect 268988 423308 268994 423360
rect 300026 423308 300032 423360
rect 300084 423348 300090 423360
rect 331214 423348 331220 423360
rect 300084 423320 331220 423348
rect 300084 423308 300090 423320
rect 331214 423308 331220 423320
rect 331272 423308 331278 423360
rect 137922 423240 137928 423292
rect 137980 423280 137986 423292
rect 313366 423280 313372 423292
rect 137980 423252 313372 423280
rect 137980 423240 137986 423252
rect 313366 423240 313372 423252
rect 313424 423240 313430 423292
rect 89622 423172 89628 423224
rect 89680 423212 89686 423224
rect 273346 423212 273352 423224
rect 89680 423184 273352 423212
rect 89680 423172 89686 423184
rect 273346 423172 273352 423184
rect 273404 423172 273410 423224
rect 295610 423172 295616 423224
rect 295668 423212 295674 423224
rect 397454 423212 397460 423224
rect 295668 423184 397460 423212
rect 295668 423172 295674 423184
rect 397454 423172 397460 423184
rect 397512 423172 397518 423224
rect 246666 423104 246672 423156
rect 246724 423144 246730 423156
rect 477494 423144 477500 423156
rect 246724 423116 477500 423144
rect 246724 423104 246730 423116
rect 477494 423104 477500 423116
rect 477552 423104 477558 423156
rect 73062 423036 73068 423088
rect 73120 423076 73126 423088
rect 317782 423076 317788 423088
rect 73120 423048 317788 423076
rect 73120 423036 73126 423048
rect 317782 423036 317788 423048
rect 317840 423036 317846 423088
rect 24762 422968 24768 423020
rect 24820 423008 24826 423020
rect 277762 423008 277768 423020
rect 24820 422980 277768 423008
rect 24820 422968 24826 422980
rect 277762 422968 277768 422980
rect 277820 422968 277826 423020
rect 286686 422968 286692 423020
rect 286744 423008 286750 423020
rect 527174 423008 527180 423020
rect 286744 422980 527180 423008
rect 286744 422968 286750 422980
rect 527174 422968 527180 422980
rect 527232 422968 527238 423020
rect 242250 422900 242256 422952
rect 242308 422940 242314 422952
rect 542354 422940 542360 422952
rect 242308 422912 542360 422940
rect 242308 422900 242314 422912
rect 542354 422900 542360 422912
rect 542412 422900 542418 422952
rect 255590 422424 255596 422476
rect 255648 422464 255654 422476
rect 256602 422464 256608 422476
rect 255648 422436 256608 422464
rect 255648 422424 255654 422436
rect 256602 422424 256608 422436
rect 256660 422424 256666 422476
rect 321830 419432 321836 419484
rect 321888 419472 321894 419484
rect 338758 419472 338764 419484
rect 321888 419444 338764 419472
rect 321888 419432 321894 419444
rect 338758 419432 338764 419444
rect 338816 419432 338822 419484
rect 321830 416712 321836 416764
rect 321888 416752 321894 416764
rect 393958 416752 393964 416764
rect 321888 416724 393964 416752
rect 321888 416712 321894 416724
rect 393958 416712 393964 416724
rect 394016 416712 394022 416764
rect 394050 415420 394056 415472
rect 394108 415460 394114 415472
rect 579614 415460 579620 415472
rect 394108 415432 579620 415460
rect 394108 415420 394114 415432
rect 579614 415420 579620 415432
rect 579672 415420 579678 415472
rect 17218 413992 17224 414044
rect 17276 414032 17282 414044
rect 237374 414032 237380 414044
rect 17276 414004 237380 414032
rect 17276 413992 17282 414004
rect 237374 413992 237380 414004
rect 237432 413992 237438 414044
rect 322198 413924 322204 413976
rect 322256 413964 322262 413976
rect 384298 413964 384304 413976
rect 322256 413936 384304 413964
rect 322256 413924 322262 413936
rect 384298 413924 384304 413936
rect 384356 413924 384362 413976
rect 322198 411204 322204 411256
rect 322256 411244 322262 411256
rect 380158 411244 380164 411256
rect 322256 411216 380164 411244
rect 322256 411204 322262 411216
rect 380158 411204 380164 411216
rect 380216 411204 380222 411256
rect 15838 408484 15844 408536
rect 15896 408524 15902 408536
rect 237374 408524 237380 408536
rect 15896 408496 237380 408524
rect 15896 408484 15902 408496
rect 237374 408484 237380 408496
rect 237432 408484 237438 408536
rect 322014 408416 322020 408468
rect 322072 408456 322078 408468
rect 395338 408456 395344 408468
rect 322072 408428 395344 408456
rect 322072 408416 322078 408428
rect 395338 408416 395344 408428
rect 395396 408416 395402 408468
rect 57238 405696 57244 405748
rect 57296 405736 57302 405748
rect 237374 405736 237380 405748
rect 57296 405708 237380 405736
rect 57296 405696 57302 405708
rect 237374 405696 237380 405708
rect 237432 405696 237438 405748
rect 321830 405628 321836 405680
rect 321888 405668 321894 405680
rect 394050 405668 394056 405680
rect 321888 405640 394056 405668
rect 321888 405628 321894 405640
rect 394050 405628 394056 405640
rect 394108 405628 394114 405680
rect 13078 402976 13084 403028
rect 13136 403016 13142 403028
rect 237374 403016 237380 403028
rect 13136 402988 237380 403016
rect 13136 402976 13142 402988
rect 237374 402976 237380 402988
rect 237432 402976 237438 403028
rect 46198 398828 46204 398880
rect 46256 398868 46262 398880
rect 237374 398868 237380 398880
rect 46256 398840 237380 398868
rect 46256 398828 46262 398840
rect 237374 398828 237380 398840
rect 237432 398828 237438 398880
rect 10410 396040 10416 396092
rect 10468 396080 10474 396092
rect 237374 396080 237380 396092
rect 10468 396052 237380 396080
rect 10468 396040 10474 396052
rect 237374 396040 237380 396052
rect 237432 396040 237438 396092
rect 322198 396040 322204 396092
rect 322256 396080 322262 396092
rect 334618 396080 334624 396092
rect 322256 396052 334624 396080
rect 322256 396040 322262 396052
rect 334618 396040 334624 396052
rect 334676 396040 334682 396092
rect 322474 394612 322480 394664
rect 322532 394652 322538 394664
rect 580258 394652 580264 394664
rect 322532 394624 580264 394652
rect 322532 394612 322538 394624
rect 580258 394612 580264 394624
rect 580316 394612 580322 394664
rect 322474 391892 322480 391944
rect 322532 391932 322538 391944
rect 580350 391932 580356 391944
rect 322532 391904 580356 391932
rect 322532 391892 322538 391904
rect 580350 391892 580356 391904
rect 580408 391892 580414 391944
rect 6178 390464 6184 390516
rect 6236 390504 6242 390516
rect 237374 390504 237380 390516
rect 6236 390476 237380 390504
rect 6236 390464 6242 390476
rect 237374 390464 237380 390476
rect 237432 390464 237438 390516
rect 322474 389104 322480 389156
rect 322532 389144 322538 389156
rect 580442 389144 580448 389156
rect 322532 389116 580448 389144
rect 322532 389104 322538 389116
rect 580442 389104 580448 389116
rect 580500 389104 580506 389156
rect 3878 387744 3884 387796
rect 3936 387784 3942 387796
rect 237374 387784 237380 387796
rect 3936 387756 237380 387784
rect 3936 387744 3942 387756
rect 237374 387744 237380 387756
rect 237432 387744 237438 387796
rect 322474 386316 322480 386368
rect 322532 386356 322538 386368
rect 391198 386356 391204 386368
rect 322532 386328 391204 386356
rect 322532 386316 322538 386328
rect 391198 386316 391204 386328
rect 391256 386316 391262 386368
rect 3786 384956 3792 385008
rect 3844 384996 3850 385008
rect 237374 384996 237380 385008
rect 3844 384968 237380 384996
rect 3844 384956 3850 384968
rect 237374 384956 237380 384968
rect 237432 384956 237438 385008
rect 322474 383596 322480 383648
rect 322532 383636 322538 383648
rect 388438 383636 388444 383648
rect 322532 383608 388444 383636
rect 322532 383596 322538 383608
rect 388438 383596 388444 383608
rect 388496 383596 388502 383648
rect 3602 382168 3608 382220
rect 3660 382208 3666 382220
rect 237374 382208 237380 382220
rect 3660 382180 237380 382208
rect 3660 382168 3666 382180
rect 237374 382168 237380 382180
rect 237432 382168 237438 382220
rect 322474 380808 322480 380860
rect 322532 380848 322538 380860
rect 580534 380848 580540 380860
rect 322532 380820 580540 380848
rect 322532 380808 322538 380820
rect 580534 380808 580540 380820
rect 580592 380808 580598 380860
rect 3510 378088 3516 378140
rect 3568 378128 3574 378140
rect 237374 378128 237380 378140
rect 3568 378100 237380 378128
rect 3568 378088 3574 378100
rect 237374 378088 237380 378100
rect 237432 378088 237438 378140
rect 322474 378088 322480 378140
rect 322532 378128 322538 378140
rect 580626 378128 580632 378140
rect 322532 378100 580632 378128
rect 322532 378088 322538 378100
rect 580626 378088 580632 378100
rect 580684 378088 580690 378140
rect 8202 375300 8208 375352
rect 8260 375340 8266 375352
rect 237374 375340 237380 375352
rect 8260 375312 237380 375340
rect 8260 375300 8266 375312
rect 237374 375300 237380 375312
rect 237432 375300 237438 375352
rect 33778 371220 33784 371272
rect 33836 371260 33842 371272
rect 237374 371260 237380 371272
rect 33836 371232 237380 371260
rect 33836 371220 33842 371232
rect 237374 371220 237380 371232
rect 237432 371220 237438 371272
rect 321830 371220 321836 371272
rect 321888 371260 321894 371272
rect 355318 371260 355324 371272
rect 321888 371232 355324 371260
rect 321888 371220 321894 371232
rect 355318 371220 355324 371232
rect 355376 371220 355382 371272
rect 322198 369792 322204 369844
rect 322256 369832 322262 369844
rect 580166 369832 580172 369844
rect 322256 369804 580172 369832
rect 322256 369792 322262 369804
rect 580166 369792 580172 369804
rect 580224 369792 580230 369844
rect 2958 367004 2964 367056
rect 3016 367044 3022 367056
rect 238294 367044 238300 367056
rect 3016 367016 238300 367044
rect 3016 367004 3022 367016
rect 238294 367004 238300 367016
rect 238352 367004 238358 367056
rect 31018 365712 31024 365764
rect 31076 365752 31082 365764
rect 237374 365752 237380 365764
rect 31076 365724 237380 365752
rect 31076 365712 31082 365724
rect 237374 365712 237380 365724
rect 237432 365712 237438 365764
rect 321830 362924 321836 362976
rect 321888 362964 321894 362976
rect 348418 362964 348424 362976
rect 321888 362936 348424 362964
rect 321888 362924 321894 362936
rect 348418 362924 348424 362936
rect 348476 362924 348482 362976
rect 321830 360204 321836 360256
rect 321888 360244 321894 360256
rect 333238 360244 333244 360256
rect 321888 360216 333244 360244
rect 321888 360204 321894 360216
rect 333238 360204 333244 360216
rect 333296 360204 333302 360256
rect 28258 358776 28264 358828
rect 28316 358816 28322 358828
rect 237374 358816 237380 358828
rect 28316 358788 237380 358816
rect 28316 358776 28322 358788
rect 237374 358776 237380 358788
rect 237432 358776 237438 358828
rect 322290 358708 322296 358760
rect 322348 358748 322354 358760
rect 579982 358748 579988 358760
rect 322348 358720 579988 358748
rect 322348 358708 322354 358720
rect 579982 358708 579988 358720
rect 580040 358708 580046 358760
rect 321646 355104 321652 355156
rect 321704 355144 321710 355156
rect 326338 355144 326344 355156
rect 321704 355116 326344 355144
rect 321704 355104 321710 355116
rect 326338 355104 326344 355116
rect 326396 355104 326402 355156
rect 6178 351908 6184 351960
rect 6236 351948 6242 351960
rect 237374 351948 237380 351960
rect 6236 351920 237380 351948
rect 6236 351908 6242 351920
rect 237374 351908 237380 351920
rect 237432 351908 237438 351960
rect 322014 349120 322020 349172
rect 322072 349160 322078 349172
rect 341518 349160 341524 349172
rect 322072 349132 341524 349160
rect 322072 349120 322078 349132
rect 341518 349120 341524 349132
rect 341576 349120 341582 349172
rect 3602 347692 3608 347744
rect 3660 347732 3666 347744
rect 237374 347732 237380 347744
rect 3660 347704 237380 347732
rect 3660 347692 3666 347704
rect 237374 347692 237380 347704
rect 237432 347692 237438 347744
rect 322014 346400 322020 346452
rect 322072 346440 322078 346452
rect 384298 346440 384304 346452
rect 322072 346412 384304 346440
rect 322072 346400 322078 346412
rect 384298 346400 384304 346412
rect 384356 346400 384362 346452
rect 322290 345040 322296 345092
rect 322348 345080 322354 345092
rect 327718 345080 327724 345092
rect 322348 345052 327724 345080
rect 322348 345040 322354 345052
rect 327718 345040 327724 345052
rect 327776 345040 327782 345092
rect 21358 344972 21364 345024
rect 21416 345012 21422 345024
rect 237374 345012 237380 345024
rect 21416 344984 237380 345012
rect 21416 344972 21422 344984
rect 237374 344972 237380 344984
rect 237432 344972 237438 345024
rect 3694 340824 3700 340876
rect 3752 340864 3758 340876
rect 237374 340864 237380 340876
rect 3752 340836 237380 340864
rect 3752 340824 3758 340836
rect 237374 340824 237380 340836
rect 237432 340824 237438 340876
rect 322290 339464 322296 339516
rect 322348 339504 322354 339516
rect 406378 339504 406384 339516
rect 322348 339476 406384 339504
rect 322348 339464 322354 339476
rect 406378 339464 406384 339476
rect 406436 339464 406442 339516
rect 19978 338036 19984 338088
rect 20036 338076 20042 338088
rect 237374 338076 237380 338088
rect 20036 338048 237380 338076
rect 20036 338036 20042 338048
rect 237374 338036 237380 338048
rect 237432 338036 237438 338088
rect 3418 335248 3424 335300
rect 3476 335288 3482 335300
rect 237374 335288 237380 335300
rect 3476 335260 237380 335288
rect 3476 335248 3482 335260
rect 237374 335248 237380 335260
rect 237432 335248 237438 335300
rect 322106 333956 322112 334008
rect 322164 333996 322170 334008
rect 340138 333996 340144 334008
rect 322164 333968 340144 333996
rect 322164 333956 322170 333968
rect 340138 333956 340144 333968
rect 340196 333956 340202 334008
rect 14458 332528 14464 332580
rect 14516 332568 14522 332580
rect 237374 332568 237380 332580
rect 14516 332540 237380 332568
rect 14516 332528 14522 332540
rect 237374 332528 237380 332540
rect 237432 332528 237438 332580
rect 322106 331236 322112 331288
rect 322164 331276 322170 331288
rect 429838 331276 429844 331288
rect 322164 331248 429844 331276
rect 322164 331236 322170 331248
rect 429838 331236 429844 331248
rect 429896 331236 429902 331288
rect 314378 328312 314384 328364
rect 314436 328352 314442 328364
rect 320910 328352 320916 328364
rect 314436 328324 320916 328352
rect 314436 328312 314442 328324
rect 320910 328312 320916 328324
rect 320968 328312 320974 328364
rect 312354 328176 312360 328228
rect 312412 328216 312418 328228
rect 323578 328216 323584 328228
rect 312412 328188 323584 328216
rect 312412 328176 312418 328188
rect 323578 328176 323584 328188
rect 323636 328176 323642 328228
rect 239398 328108 239404 328160
rect 239456 328148 239462 328160
rect 254118 328148 254124 328160
rect 239456 328120 254124 328148
rect 239456 328108 239462 328120
rect 254118 328108 254124 328120
rect 254176 328108 254182 328160
rect 279421 328151 279479 328157
rect 279421 328117 279433 328151
rect 279467 328148 279479 328151
rect 285858 328148 285864 328160
rect 279467 328120 285864 328148
rect 279467 328117 279479 328120
rect 279421 328111 279479 328117
rect 285858 328108 285864 328120
rect 285916 328108 285922 328160
rect 302602 328108 302608 328160
rect 302660 328148 302666 328160
rect 312538 328148 312544 328160
rect 302660 328120 312544 328148
rect 302660 328108 302666 328120
rect 312538 328108 312544 328120
rect 312596 328108 312602 328160
rect 229738 328040 229744 328092
rect 229796 328080 229802 328092
rect 246390 328080 246396 328092
rect 229796 328052 246396 328080
rect 229796 328040 229802 328052
rect 246390 328040 246396 328052
rect 246448 328040 246454 328092
rect 249061 328083 249119 328089
rect 249061 328049 249073 328083
rect 249107 328080 249119 328083
rect 254486 328080 254492 328092
rect 249107 328052 254492 328080
rect 249107 328049 249119 328052
rect 249061 328043 249119 328049
rect 254486 328040 254492 328052
rect 254544 328040 254550 328092
rect 272518 328040 272524 328092
rect 272576 328080 272582 328092
rect 280798 328080 280804 328092
rect 272576 328052 280804 328080
rect 272576 328040 272582 328052
rect 280798 328040 280804 328052
rect 280856 328040 280862 328092
rect 307018 328040 307024 328092
rect 307076 328080 307082 328092
rect 315853 328083 315911 328089
rect 315853 328080 315865 328083
rect 307076 328052 315865 328080
rect 307076 328040 307082 328052
rect 315853 328049 315865 328052
rect 315899 328049 315911 328083
rect 315853 328043 315911 328049
rect 236638 327972 236644 328024
rect 236696 328012 236702 328024
rect 258534 328012 258540 328024
rect 236696 327984 258540 328012
rect 236696 327972 236702 327984
rect 258534 327972 258540 327984
rect 258592 327972 258598 328024
rect 277394 327972 277400 328024
rect 277452 328012 277458 328024
rect 277670 328012 277676 328024
rect 277452 327984 277676 328012
rect 277452 327972 277458 327984
rect 277670 327972 277676 327984
rect 277728 327972 277734 328024
rect 279510 327972 279516 328024
rect 279568 328012 279574 328024
rect 289078 328012 289084 328024
rect 279568 327984 289084 328012
rect 279568 327972 279574 327984
rect 289078 327972 289084 327984
rect 289136 327972 289142 328024
rect 293954 327972 293960 328024
rect 294012 328012 294018 328024
rect 294322 328012 294328 328024
rect 294012 327984 294328 328012
rect 294012 327972 294018 327984
rect 294322 327972 294328 327984
rect 294380 327972 294386 328024
rect 300946 327972 300952 328024
rect 301004 328012 301010 328024
rect 301866 328012 301872 328024
rect 301004 327984 301872 328012
rect 301004 327972 301010 327984
rect 301866 327972 301872 327984
rect 301924 327972 301930 328024
rect 306190 327972 306196 328024
rect 306248 328012 306254 328024
rect 345014 328012 345020 328024
rect 306248 327984 345020 328012
rect 306248 327972 306254 327984
rect 345014 327972 345020 327984
rect 345072 327972 345078 328024
rect 231118 327904 231124 327956
rect 231176 327944 231182 327956
rect 249061 327947 249119 327953
rect 249061 327944 249073 327947
rect 231176 327916 249073 327944
rect 231176 327904 231182 327916
rect 249061 327913 249073 327916
rect 249107 327913 249119 327947
rect 249061 327907 249119 327913
rect 258718 327904 258724 327956
rect 258776 327944 258782 327956
rect 267918 327944 267924 327956
rect 258776 327916 267924 327944
rect 258776 327904 258782 327916
rect 267918 327904 267924 327916
rect 267976 327904 267982 327956
rect 272058 327904 272064 327956
rect 272116 327944 272122 327956
rect 273162 327944 273168 327956
rect 272116 327916 273168 327944
rect 272116 327904 272122 327916
rect 273162 327904 273168 327916
rect 273220 327904 273226 327956
rect 276934 327904 276940 327956
rect 276992 327944 276998 327956
rect 317509 327947 317567 327953
rect 317509 327944 317521 327947
rect 276992 327916 317521 327944
rect 276992 327904 276998 327916
rect 317509 327913 317521 327916
rect 317555 327913 317567 327947
rect 317509 327907 317567 327913
rect 317598 327904 317604 327956
rect 317656 327944 317662 327956
rect 318426 327944 318432 327956
rect 317656 327916 318432 327944
rect 317656 327904 317662 327916
rect 318426 327904 318432 327916
rect 318484 327904 318490 327956
rect 233878 327836 233884 327888
rect 233936 327876 233942 327888
rect 259454 327876 259460 327888
rect 233936 327848 259460 327876
rect 233936 327836 233942 327848
rect 259454 327836 259460 327848
rect 259512 327836 259518 327888
rect 272886 327836 272892 327888
rect 272944 327876 272950 327888
rect 273070 327876 273076 327888
rect 272944 327848 273076 327876
rect 272944 327836 272950 327848
rect 273070 327836 273076 327848
rect 273128 327836 273134 327888
rect 273180 327848 279556 327876
rect 232498 327768 232504 327820
rect 232556 327808 232562 327820
rect 260834 327808 260840 327820
rect 232556 327780 260840 327808
rect 232556 327768 232562 327780
rect 260834 327768 260840 327780
rect 260892 327768 260898 327820
rect 268930 327768 268936 327820
rect 268988 327808 268994 327820
rect 273180 327808 273208 327848
rect 268988 327780 273208 327808
rect 268988 327768 268994 327780
rect 276658 327768 276664 327820
rect 276716 327808 276722 327820
rect 279421 327811 279479 327817
rect 279421 327808 279433 327811
rect 276716 327780 279433 327808
rect 276716 327768 276722 327780
rect 279421 327777 279433 327780
rect 279467 327777 279479 327811
rect 279528 327808 279556 327848
rect 279786 327836 279792 327888
rect 279844 327876 279850 327888
rect 280062 327876 280068 327888
rect 279844 327848 280068 327876
rect 279844 327836 279850 327848
rect 280062 327836 280068 327848
rect 280120 327836 280126 327888
rect 281718 327836 281724 327888
rect 281776 327876 281782 327888
rect 282546 327876 282552 327888
rect 281776 327848 282552 327876
rect 281776 327836 281782 327848
rect 282546 327836 282552 327848
rect 282604 327836 282610 327888
rect 283006 327836 283012 327888
rect 283064 327876 283070 327888
rect 283374 327876 283380 327888
rect 283064 327848 283380 327876
rect 283064 327836 283070 327848
rect 283374 327836 283380 327848
rect 283432 327836 283438 327888
rect 284938 327836 284944 327888
rect 284996 327876 285002 327888
rect 285766 327876 285772 327888
rect 284996 327848 285772 327876
rect 284996 327836 285002 327848
rect 285766 327836 285772 327848
rect 285824 327836 285830 327888
rect 287790 327836 287796 327888
rect 287848 327876 287854 327888
rect 288434 327876 288440 327888
rect 287848 327848 288440 327876
rect 287848 327836 287854 327848
rect 288434 327836 288440 327848
rect 288492 327836 288498 327888
rect 290458 327836 290464 327888
rect 290516 327876 290522 327888
rect 291194 327876 291200 327888
rect 290516 327848 291200 327876
rect 290516 327836 290522 327848
rect 291194 327836 291200 327848
rect 291252 327836 291258 327888
rect 291930 327836 291936 327888
rect 291988 327876 291994 327888
rect 292666 327876 292672 327888
rect 291988 327848 292672 327876
rect 291988 327836 291994 327848
rect 292666 327836 292672 327848
rect 292724 327836 292730 327888
rect 295518 327836 295524 327888
rect 295576 327876 295582 327888
rect 296346 327876 296352 327888
rect 295576 327848 296352 327876
rect 295576 327836 295582 327848
rect 296346 327836 296352 327848
rect 296404 327836 296410 327888
rect 298094 327836 298100 327888
rect 298152 327876 298158 327888
rect 298370 327876 298376 327888
rect 298152 327848 298376 327876
rect 298152 327836 298158 327848
rect 298370 327836 298376 327848
rect 298428 327836 298434 327888
rect 315206 327836 315212 327888
rect 315264 327876 315270 327888
rect 315758 327876 315764 327888
rect 315264 327848 315764 327876
rect 315264 327836 315270 327848
rect 315758 327836 315764 327848
rect 315816 327836 315822 327888
rect 315853 327879 315911 327885
rect 315853 327845 315865 327879
rect 315899 327876 315911 327879
rect 351914 327876 351920 327888
rect 315899 327848 351920 327876
rect 315899 327845 315911 327848
rect 315853 327839 315911 327845
rect 351914 327836 351920 327848
rect 351972 327836 351978 327888
rect 281534 327808 281540 327820
rect 279528 327780 281540 327808
rect 279421 327771 279479 327777
rect 281534 327768 281540 327780
rect 281592 327768 281598 327820
rect 282914 327768 282920 327820
rect 282972 327808 282978 327820
rect 283742 327808 283748 327820
rect 282972 327780 283748 327808
rect 282972 327768 282978 327780
rect 283742 327768 283748 327780
rect 283800 327768 283806 327820
rect 289906 327768 289912 327820
rect 289964 327808 289970 327820
rect 290734 327808 290740 327820
rect 289964 327780 290740 327808
rect 289964 327768 289970 327780
rect 290734 327768 290740 327780
rect 290792 327768 290798 327820
rect 307478 327768 307484 327820
rect 307536 327808 307542 327820
rect 469214 327808 469220 327820
rect 307536 327780 469220 327808
rect 307536 327768 307542 327780
rect 469214 327768 469220 327780
rect 469272 327768 469278 327820
rect 122742 327700 122748 327752
rect 122800 327740 122806 327752
rect 240686 327740 240692 327752
rect 122800 327712 240692 327740
rect 122800 327700 122806 327712
rect 240686 327700 240692 327712
rect 240744 327700 240750 327752
rect 281810 327740 281816 327752
rect 267706 327712 281816 327740
rect 262858 327632 262864 327684
rect 262916 327672 262922 327684
rect 266354 327672 266360 327684
rect 262916 327644 266360 327672
rect 262916 327632 262922 327644
rect 266354 327632 266360 327644
rect 266412 327632 266418 327684
rect 258810 327564 258816 327616
rect 258868 327604 258874 327616
rect 267706 327604 267734 327712
rect 281810 327700 281816 327712
rect 281868 327700 281874 327752
rect 285766 327700 285772 327752
rect 285824 327740 285830 327752
rect 286594 327740 286600 327752
rect 285824 327712 286600 327740
rect 285824 327700 285830 327712
rect 286594 327700 286600 327712
rect 286652 327700 286658 327752
rect 292666 327700 292672 327752
rect 292724 327740 292730 327752
rect 293126 327740 293132 327752
rect 292724 327712 293132 327740
rect 292724 327700 292730 327712
rect 293126 327700 293132 327712
rect 293184 327700 293190 327752
rect 299566 327700 299572 327752
rect 299624 327740 299630 327752
rect 300026 327740 300032 327752
rect 299624 327712 300032 327740
rect 299624 327700 299630 327712
rect 300026 327700 300032 327712
rect 300084 327700 300090 327752
rect 302970 327700 302976 327752
rect 303028 327740 303034 327752
rect 303430 327740 303436 327752
rect 303028 327712 303436 327740
rect 303028 327700 303034 327712
rect 303430 327700 303436 327712
rect 303488 327700 303494 327752
rect 308214 327700 308220 327752
rect 308272 327740 308278 327752
rect 477494 327740 477500 327752
rect 308272 327712 477500 327740
rect 308272 327700 308278 327712
rect 477494 327700 477500 327712
rect 477552 327700 477558 327752
rect 271322 327632 271328 327684
rect 271380 327672 271386 327684
rect 271782 327672 271788 327684
rect 271380 327644 271788 327672
rect 271380 327632 271386 327644
rect 271782 327632 271788 327644
rect 271840 327632 271846 327684
rect 274082 327632 274088 327684
rect 274140 327672 274146 327684
rect 274542 327672 274548 327684
rect 274140 327644 274548 327672
rect 274140 327632 274146 327644
rect 274542 327632 274548 327644
rect 274600 327632 274606 327684
rect 278958 327632 278964 327684
rect 279016 327672 279022 327684
rect 279786 327672 279792 327684
rect 279016 327644 279792 327672
rect 279016 327632 279022 327644
rect 279786 327632 279792 327644
rect 279844 327632 279850 327684
rect 287698 327632 287704 327684
rect 287756 327672 287762 327684
rect 288618 327672 288624 327684
rect 287756 327644 288624 327672
rect 287756 327632 287762 327644
rect 288618 327632 288624 327644
rect 288676 327632 288682 327684
rect 294598 327632 294604 327684
rect 294656 327672 294662 327684
rect 295610 327672 295616 327684
rect 294656 327644 295616 327672
rect 294656 327632 294662 327644
rect 295610 327632 295616 327644
rect 295668 327632 295674 327684
rect 316402 327632 316408 327684
rect 316460 327672 316466 327684
rect 317138 327672 317144 327684
rect 316460 327644 317144 327672
rect 316460 327632 316466 327644
rect 317138 327632 317144 327644
rect 317196 327632 317202 327684
rect 317966 327632 317972 327684
rect 318024 327672 318030 327684
rect 318518 327672 318524 327684
rect 318024 327644 318524 327672
rect 318024 327632 318030 327644
rect 318518 327632 318524 327644
rect 318576 327632 318582 327684
rect 319254 327632 319260 327684
rect 319312 327672 319318 327684
rect 319898 327672 319904 327684
rect 319312 327644 319904 327672
rect 319312 327632 319318 327644
rect 319898 327632 319904 327644
rect 319956 327632 319962 327684
rect 258868 327576 267734 327604
rect 258868 327564 258874 327576
rect 291838 327564 291844 327616
rect 291896 327604 291902 327616
rect 295334 327604 295340 327616
rect 291896 327576 295340 327604
rect 291896 327564 291902 327576
rect 295334 327564 295340 327576
rect 295392 327564 295398 327616
rect 304166 327564 304172 327616
rect 304224 327604 304230 327616
rect 304810 327604 304816 327616
rect 304224 327576 304816 327604
rect 304224 327564 304230 327576
rect 304810 327564 304816 327576
rect 304868 327564 304874 327616
rect 317509 327607 317567 327613
rect 317509 327573 317521 327607
rect 317555 327604 317567 327607
rect 320818 327604 320824 327616
rect 317555 327576 320824 327604
rect 317555 327573 317567 327576
rect 317509 327567 317567 327573
rect 320818 327564 320824 327576
rect 320876 327564 320882 327616
rect 262030 327496 262036 327548
rect 262088 327536 262094 327548
rect 263594 327536 263600 327548
rect 262088 327508 263600 327536
rect 262088 327496 262094 327508
rect 263594 327496 263600 327508
rect 263652 327496 263658 327548
rect 273714 327496 273720 327548
rect 273772 327536 273778 327548
rect 274450 327536 274456 327548
rect 273772 327508 274456 327536
rect 273772 327496 273778 327508
rect 274450 327496 274456 327508
rect 274508 327496 274514 327548
rect 279418 327496 279424 327548
rect 279476 327536 279482 327548
rect 279878 327536 279884 327548
rect 279476 327508 279884 327536
rect 279476 327496 279482 327508
rect 279878 327496 279884 327508
rect 279936 327496 279942 327548
rect 301314 327496 301320 327548
rect 301372 327536 301378 327548
rect 302050 327536 302056 327548
rect 301372 327508 302056 327536
rect 301372 327496 301378 327508
rect 302050 327496 302056 327508
rect 302108 327496 302114 327548
rect 304626 327496 304632 327548
rect 304684 327536 304690 327548
rect 304902 327536 304908 327548
rect 304684 327508 304908 327536
rect 304684 327496 304690 327508
rect 304902 327496 304908 327508
rect 304960 327496 304966 327548
rect 308674 327496 308680 327548
rect 308732 327536 308738 327548
rect 309042 327536 309048 327548
rect 308732 327508 309048 327536
rect 308732 327496 308738 327508
rect 309042 327496 309048 327508
rect 309100 327496 309106 327548
rect 311434 327496 311440 327548
rect 311492 327536 311498 327548
rect 311710 327536 311716 327548
rect 311492 327508 311716 327536
rect 311492 327496 311498 327508
rect 311710 327496 311716 327508
rect 311768 327496 311774 327548
rect 316770 327496 316776 327548
rect 316828 327536 316834 327548
rect 317322 327536 317328 327548
rect 316828 327508 317328 327536
rect 316828 327496 316834 327508
rect 317322 327496 317328 327508
rect 317380 327496 317386 327548
rect 315574 327428 315580 327480
rect 315632 327468 315638 327480
rect 315942 327468 315948 327480
rect 315632 327440 315948 327468
rect 315632 327428 315638 327440
rect 315942 327428 315948 327440
rect 316000 327428 316006 327480
rect 262950 327360 262956 327412
rect 263008 327400 263014 327412
rect 263870 327400 263876 327412
rect 263008 327372 263876 327400
rect 263008 327360 263014 327372
rect 263870 327360 263876 327372
rect 263928 327360 263934 327412
rect 276566 327360 276572 327412
rect 276624 327400 276630 327412
rect 277302 327400 277308 327412
rect 276624 327372 277308 327400
rect 276624 327360 276630 327372
rect 277302 327360 277308 327372
rect 277360 327360 277366 327412
rect 280614 327360 280620 327412
rect 280672 327400 280678 327412
rect 281258 327400 281264 327412
rect 280672 327372 281264 327400
rect 280672 327360 280678 327372
rect 281258 327360 281264 327372
rect 281316 327360 281322 327412
rect 305454 327360 305460 327412
rect 305512 327400 305518 327412
rect 306282 327400 306288 327412
rect 305512 327372 306288 327400
rect 305512 327360 305518 327372
rect 306282 327360 306288 327372
rect 306340 327360 306346 327412
rect 306650 327360 306656 327412
rect 306708 327400 306714 327412
rect 307570 327400 307576 327412
rect 306708 327372 307576 327400
rect 306708 327360 306714 327372
rect 307570 327360 307576 327372
rect 307628 327360 307634 327412
rect 311066 327360 311072 327412
rect 311124 327400 311130 327412
rect 311618 327400 311624 327412
rect 311124 327372 311624 327400
rect 311124 327360 311130 327372
rect 311618 327360 311624 327372
rect 311676 327360 311682 327412
rect 261938 327292 261944 327344
rect 261996 327332 262002 327344
rect 269114 327332 269120 327344
rect 261996 327304 269120 327332
rect 261996 327292 262002 327304
rect 269114 327292 269120 327304
rect 269172 327292 269178 327344
rect 279418 327292 279424 327344
rect 279476 327332 279482 327344
rect 285030 327332 285036 327344
rect 279476 327304 285036 327332
rect 279476 327292 279482 327304
rect 285030 327292 285036 327304
rect 285088 327292 285094 327344
rect 256234 327088 256240 327140
rect 256292 327128 256298 327140
rect 256694 327128 256700 327140
rect 256292 327100 256700 327128
rect 256292 327088 256298 327100
rect 256694 327088 256700 327100
rect 256752 327088 256758 327140
rect 258350 327088 258356 327140
rect 258408 327128 258414 327140
rect 259822 327128 259828 327140
rect 258408 327100 259828 327128
rect 258408 327088 258414 327100
rect 259822 327088 259828 327100
rect 259880 327088 259886 327140
rect 265618 327088 265624 327140
rect 265676 327128 265682 327140
rect 267734 327128 267740 327140
rect 265676 327100 267740 327128
rect 265676 327088 265682 327100
rect 267734 327088 267740 327100
rect 267792 327088 267798 327140
rect 268378 327088 268384 327140
rect 268436 327128 268442 327140
rect 268930 327128 268936 327140
rect 268436 327100 268936 327128
rect 268436 327088 268442 327100
rect 268930 327088 268936 327100
rect 268988 327088 268994 327140
rect 286318 327088 286324 327140
rect 286376 327128 286382 327140
rect 287146 327128 287152 327140
rect 286376 327100 287152 327128
rect 286376 327088 286382 327100
rect 287146 327088 287152 327100
rect 287204 327088 287210 327140
rect 219342 326408 219348 326460
rect 219400 326448 219406 326460
rect 264974 326448 264980 326460
rect 219400 326420 264980 326448
rect 219400 326408 219406 326420
rect 264974 326408 264980 326420
rect 265032 326408 265038 326460
rect 126882 326340 126888 326392
rect 126940 326380 126946 326392
rect 239398 326380 239404 326392
rect 126940 326352 239404 326380
rect 126940 326340 126946 326352
rect 239398 326340 239404 326352
rect 239456 326340 239462 326392
rect 274910 326340 274916 326392
rect 274968 326380 274974 326392
rect 305086 326380 305092 326392
rect 274968 326352 305092 326380
rect 274968 326340 274974 326352
rect 305086 326340 305092 326352
rect 305144 326340 305150 326392
rect 309318 326340 309324 326392
rect 309376 326380 309382 326392
rect 487154 326380 487160 326392
rect 309376 326352 487160 326380
rect 309376 326340 309382 326352
rect 487154 326340 487160 326352
rect 487212 326340 487218 326392
rect 262398 326272 262404 326324
rect 262456 326272 262462 326324
rect 262416 326108 262444 326272
rect 262490 326108 262496 326120
rect 262416 326080 262496 326108
rect 262490 326068 262496 326080
rect 262548 326068 262554 326120
rect 247310 325864 247316 325916
rect 247368 325864 247374 325916
rect 248598 325904 248604 325916
rect 248559 325876 248604 325904
rect 248598 325864 248604 325876
rect 248656 325864 248662 325916
rect 240410 325728 240416 325780
rect 240468 325768 240474 325780
rect 241054 325768 241060 325780
rect 240468 325740 241060 325768
rect 240468 325728 240474 325740
rect 241054 325728 241060 325740
rect 241112 325728 241118 325780
rect 241514 325728 241520 325780
rect 241572 325768 241578 325780
rect 242342 325768 242348 325780
rect 241572 325740 242348 325768
rect 241572 325728 241578 325740
rect 242342 325728 242348 325740
rect 242400 325728 242406 325780
rect 244366 325728 244372 325780
rect 244424 325768 244430 325780
rect 244734 325768 244740 325780
rect 244424 325740 244740 325768
rect 244424 325728 244430 325740
rect 244734 325728 244740 325740
rect 244792 325728 244798 325780
rect 247328 325712 247356 325864
rect 247586 325728 247592 325780
rect 247644 325768 247650 325780
rect 248046 325768 248052 325780
rect 247644 325740 248052 325768
rect 247644 325728 247650 325740
rect 248046 325728 248052 325740
rect 248104 325728 248110 325780
rect 248414 325728 248420 325780
rect 248472 325768 248478 325780
rect 249242 325768 249248 325780
rect 248472 325740 249248 325768
rect 248472 325728 248478 325740
rect 249242 325728 249248 325740
rect 249300 325728 249306 325780
rect 251634 325728 251640 325780
rect 251692 325768 251698 325780
rect 252094 325768 252100 325780
rect 251692 325740 252100 325768
rect 251692 325728 251698 325740
rect 252094 325728 252100 325740
rect 252152 325728 252158 325780
rect 252554 325728 252560 325780
rect 252612 325768 252618 325780
rect 253290 325768 253296 325780
rect 252612 325740 253296 325768
rect 252612 325728 252618 325740
rect 253290 325728 253296 325740
rect 253348 325728 253354 325780
rect 247310 325660 247316 325712
rect 247368 325660 247374 325712
rect 262306 325660 262312 325712
rect 262364 325700 262370 325712
rect 263042 325700 263048 325712
rect 262364 325672 263048 325700
rect 262364 325660 262370 325672
rect 263042 325660 263048 325672
rect 263100 325660 263106 325712
rect 243354 325632 243360 325644
rect 243280 325604 243360 325632
rect 243280 325440 243308 325604
rect 243354 325592 243360 325604
rect 243412 325592 243418 325644
rect 257154 325632 257160 325644
rect 257080 325604 257160 325632
rect 257080 325440 257108 325604
rect 257154 325592 257160 325604
rect 257212 325592 257218 325644
rect 243262 325388 243268 325440
rect 243320 325388 243326 325440
rect 257062 325388 257068 325440
rect 257120 325388 257126 325440
rect 162762 324912 162768 324964
rect 162820 324952 162826 324964
rect 258258 324952 258264 324964
rect 162820 324924 258264 324952
rect 162820 324912 162826 324924
rect 258258 324912 258264 324924
rect 258316 324912 258322 324964
rect 275002 324912 275008 324964
rect 275060 324952 275066 324964
rect 307754 324952 307760 324964
rect 275060 324924 307760 324952
rect 275060 324912 275066 324924
rect 307754 324912 307760 324924
rect 307812 324912 307818 324964
rect 309410 324912 309416 324964
rect 309468 324952 309474 324964
rect 491294 324952 491300 324964
rect 309468 324924 491300 324952
rect 309468 324912 309474 324924
rect 491294 324912 491300 324924
rect 491352 324912 491358 324964
rect 3234 324232 3240 324284
rect 3292 324272 3298 324284
rect 238478 324272 238484 324284
rect 3292 324244 238484 324272
rect 3292 324232 3298 324244
rect 238478 324232 238484 324244
rect 238536 324232 238542 324284
rect 243170 323620 243176 323672
rect 243228 323660 243234 323672
rect 243538 323660 243544 323672
rect 243228 323632 243544 323660
rect 243228 323620 243234 323632
rect 243538 323620 243544 323632
rect 243596 323620 243602 323672
rect 247218 323620 247224 323672
rect 247276 323660 247282 323672
rect 247402 323660 247408 323672
rect 247276 323632 247408 323660
rect 247276 323620 247282 323632
rect 247402 323620 247408 323632
rect 247460 323620 247466 323672
rect 248598 323660 248604 323672
rect 248559 323632 248604 323660
rect 248598 323620 248604 323632
rect 248656 323620 248662 323672
rect 277486 323620 277492 323672
rect 277544 323660 277550 323672
rect 329834 323660 329840 323672
rect 277544 323632 329840 323660
rect 277544 323620 277550 323632
rect 329834 323620 329840 323632
rect 329892 323620 329898 323672
rect 227622 323552 227628 323604
rect 227680 323592 227686 323604
rect 265158 323592 265164 323604
rect 227680 323564 265164 323592
rect 227680 323552 227686 323564
rect 265158 323552 265164 323564
rect 265216 323552 265222 323604
rect 310606 323552 310612 323604
rect 310664 323592 310670 323604
rect 498194 323592 498200 323604
rect 310664 323564 498200 323592
rect 310664 323552 310670 323564
rect 498194 323552 498200 323564
rect 498252 323552 498258 323604
rect 322750 322872 322756 322924
rect 322808 322912 322814 322924
rect 580166 322912 580172 322924
rect 322808 322884 580172 322912
rect 322808 322872 322814 322884
rect 580166 322872 580172 322884
rect 580224 322872 580230 322924
rect 231762 322260 231768 322312
rect 231820 322300 231826 322312
rect 292758 322300 292764 322312
rect 231820 322272 292764 322300
rect 231820 322260 231826 322272
rect 292758 322260 292764 322272
rect 292816 322260 292822 322312
rect 169662 322192 169668 322244
rect 169720 322232 169726 322244
rect 258994 322232 259000 322244
rect 169720 322204 259000 322232
rect 169720 322192 169726 322204
rect 258994 322192 259000 322204
rect 259052 322192 259058 322244
rect 300946 322192 300952 322244
rect 301004 322232 301010 322244
rect 309134 322232 309140 322244
rect 301004 322204 309140 322232
rect 301004 322192 301010 322204
rect 309134 322192 309140 322204
rect 309192 322192 309198 322244
rect 277394 320900 277400 320952
rect 277452 320940 277458 320952
rect 332594 320940 332600 320952
rect 277452 320912 332600 320940
rect 277452 320900 277458 320912
rect 332594 320900 332600 320912
rect 332652 320900 332658 320952
rect 176562 320832 176568 320884
rect 176620 320872 176626 320884
rect 258350 320872 258356 320884
rect 176620 320844 258356 320872
rect 176620 320832 176626 320844
rect 258350 320832 258356 320844
rect 258408 320832 258414 320884
rect 313366 320832 313372 320884
rect 313424 320872 313430 320884
rect 523034 320872 523040 320884
rect 313424 320844 523040 320872
rect 313424 320832 313430 320844
rect 523034 320832 523040 320844
rect 523092 320832 523098 320884
rect 278038 319472 278044 319524
rect 278096 319512 278102 319524
rect 336734 319512 336740 319524
rect 278096 319484 336740 319512
rect 278096 319472 278102 319484
rect 336734 319472 336740 319484
rect 336792 319472 336798 319524
rect 180702 319404 180708 319456
rect 180760 319444 180766 319456
rect 260190 319444 260196 319456
rect 180760 319416 260196 319444
rect 180760 319404 180766 319416
rect 260190 319404 260196 319416
rect 260248 319404 260254 319456
rect 313550 319404 313556 319456
rect 313608 319444 313614 319456
rect 527174 319444 527180 319456
rect 313608 319416 527180 319444
rect 313608 319404 313614 319416
rect 527174 319404 527180 319416
rect 527232 319404 527238 319456
rect 262214 318996 262220 319048
rect 262272 319036 262278 319048
rect 262582 319036 262588 319048
rect 262272 319008 262588 319036
rect 262272 318996 262278 319008
rect 262582 318996 262588 319008
rect 262640 318996 262646 319048
rect 256970 318792 256976 318844
rect 257028 318832 257034 318844
rect 257338 318832 257344 318844
rect 257028 318804 257344 318832
rect 257028 318792 257034 318804
rect 257338 318792 257344 318804
rect 257396 318792 257402 318844
rect 279786 318112 279792 318164
rect 279844 318152 279850 318164
rect 339494 318152 339500 318164
rect 279844 318124 339500 318152
rect 279844 318112 279850 318124
rect 339494 318112 339500 318124
rect 339552 318112 339558 318164
rect 187602 318044 187608 318096
rect 187660 318084 187666 318096
rect 261018 318084 261024 318096
rect 187660 318056 261024 318084
rect 187660 318044 187666 318056
rect 261018 318044 261024 318056
rect 261076 318044 261082 318096
rect 318426 318044 318432 318096
rect 318484 318084 318490 318096
rect 558178 318084 558184 318096
rect 318484 318056 558184 318084
rect 318484 318044 318490 318056
rect 558178 318044 558184 318056
rect 558236 318044 558242 318096
rect 279878 316752 279884 316804
rect 279936 316792 279942 316804
rect 343634 316792 343640 316804
rect 279936 316764 343640 316792
rect 279936 316752 279942 316764
rect 343634 316752 343640 316764
rect 343692 316752 343698 316804
rect 194502 316684 194508 316736
rect 194560 316724 194566 316736
rect 261386 316724 261392 316736
rect 194560 316696 261392 316724
rect 194560 316684 194566 316696
rect 261386 316684 261392 316696
rect 261444 316684 261450 316736
rect 318518 316684 318524 316736
rect 318576 316724 318582 316736
rect 563054 316724 563060 316736
rect 318576 316696 563060 316724
rect 318576 316684 318582 316696
rect 563054 316684 563060 316696
rect 563112 316684 563118 316736
rect 198642 315256 198648 315308
rect 198700 315296 198706 315308
rect 262398 315296 262404 315308
rect 198700 315268 262404 315296
rect 198700 315256 198706 315268
rect 262398 315256 262404 315268
rect 262456 315256 262462 315308
rect 279970 315256 279976 315308
rect 280028 315296 280034 315308
rect 350534 315296 350540 315308
rect 280028 315268 350540 315296
rect 280028 315256 280034 315268
rect 350534 315256 350540 315268
rect 350592 315256 350598 315308
rect 205542 313964 205548 314016
rect 205600 314004 205606 314016
rect 262306 314004 262312 314016
rect 205600 313976 262312 314004
rect 205600 313964 205606 313976
rect 262306 313964 262312 313976
rect 262364 313964 262370 314016
rect 104802 313896 104808 313948
rect 104860 313936 104866 313948
rect 244274 313936 244280 313948
rect 104860 313908 244280 313936
rect 104860 313896 104866 313908
rect 244274 313896 244280 313908
rect 244332 313896 244338 313948
rect 311618 313896 311624 313948
rect 311676 313936 311682 313948
rect 502334 313936 502340 313948
rect 311676 313908 502340 313936
rect 311676 313896 311682 313908
rect 502334 313896 502340 313908
rect 502392 313896 502398 313948
rect 209682 312604 209688 312656
rect 209740 312644 209746 312656
rect 261570 312644 261576 312656
rect 209740 312616 261576 312644
rect 209740 312604 209746 312616
rect 261570 312604 261576 312616
rect 261628 312604 261634 312656
rect 86862 312536 86868 312588
rect 86920 312576 86926 312588
rect 241882 312576 241888 312588
rect 86920 312548 241888 312576
rect 86920 312536 86926 312548
rect 241882 312536 241888 312548
rect 241940 312536 241946 312588
rect 260742 312536 260748 312588
rect 260800 312576 260806 312588
rect 295702 312576 295708 312588
rect 260800 312548 295708 312576
rect 260800 312536 260806 312548
rect 295702 312536 295708 312548
rect 295760 312536 295766 312588
rect 311710 312536 311716 312588
rect 311768 312576 311774 312588
rect 505094 312576 505100 312588
rect 311768 312548 505100 312576
rect 311768 312536 311774 312548
rect 505094 312536 505100 312548
rect 505152 312536 505158 312588
rect 355318 311788 355324 311840
rect 355376 311828 355382 311840
rect 580166 311828 580172 311840
rect 355376 311800 580172 311828
rect 355376 311788 355382 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 212442 311176 212448 311228
rect 212500 311216 212506 311228
rect 262950 311216 262956 311228
rect 212500 311188 262956 311216
rect 212500 311176 212506 311188
rect 262950 311176 262956 311188
rect 263008 311176 263014 311228
rect 57882 311108 57888 311160
rect 57940 311148 57946 311160
rect 247310 311148 247316 311160
rect 57940 311120 247316 311148
rect 57940 311108 57946 311120
rect 247310 311108 247316 311120
rect 247368 311108 247374 311160
rect 216582 309816 216588 309868
rect 216640 309856 216646 309868
rect 263870 309856 263876 309868
rect 216640 309828 263876 309856
rect 216640 309816 216646 309828
rect 263870 309816 263876 309828
rect 263928 309816 263934 309868
rect 50982 309748 50988 309800
rect 51040 309788 51046 309800
rect 245930 309788 245936 309800
rect 51040 309760 245936 309788
rect 51040 309748 51046 309760
rect 245930 309748 245936 309760
rect 245988 309748 245994 309800
rect 311526 309748 311532 309800
rect 311584 309788 311590 309800
rect 509234 309788 509240 309800
rect 311584 309760 509240 309788
rect 311584 309748 311590 309760
rect 509234 309748 509240 309760
rect 509292 309748 509298 309800
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 10410 309108 10416 309120
rect 3384 309080 10416 309108
rect 3384 309068 3390 309080
rect 10410 309068 10416 309080
rect 10468 309068 10474 309120
rect 223482 308456 223488 308508
rect 223540 308496 223546 308508
rect 265066 308496 265072 308508
rect 223540 308468 265072 308496
rect 223540 308456 223546 308468
rect 265066 308456 265072 308468
rect 265124 308456 265130 308508
rect 10318 308388 10324 308440
rect 10376 308428 10382 308440
rect 241606 308428 241612 308440
rect 10376 308400 241612 308428
rect 10376 308388 10382 308400
rect 241606 308388 241612 308400
rect 241664 308388 241670 308440
rect 313090 308388 313096 308440
rect 313148 308428 313154 308440
rect 516134 308428 516140 308440
rect 313148 308400 516140 308428
rect 313148 308388 313154 308400
rect 516134 308388 516140 308400
rect 516192 308388 516198 308440
rect 133782 307028 133788 307080
rect 133840 307068 133846 307080
rect 254486 307068 254492 307080
rect 133840 307040 254492 307068
rect 133840 307028 133846 307040
rect 254486 307028 254492 307040
rect 254544 307028 254550 307080
rect 314562 307028 314568 307080
rect 314620 307068 314626 307080
rect 534074 307068 534080 307080
rect 314620 307040 534080 307068
rect 314620 307028 314626 307040
rect 534074 307028 534080 307040
rect 534132 307028 534138 307080
rect 142062 305600 142068 305652
rect 142120 305640 142126 305652
rect 255406 305640 255412 305652
rect 142120 305612 255412 305640
rect 142120 305600 142126 305612
rect 255406 305600 255412 305612
rect 255464 305600 255470 305652
rect 315758 305600 315764 305652
rect 315816 305640 315822 305652
rect 536834 305640 536840 305652
rect 315816 305612 536840 305640
rect 315816 305600 315822 305612
rect 536834 305600 536840 305612
rect 536892 305600 536898 305652
rect 144822 304240 144828 304292
rect 144880 304280 144886 304292
rect 255682 304280 255688 304292
rect 144880 304252 255688 304280
rect 144880 304240 144886 304252
rect 255682 304240 255688 304252
rect 255740 304240 255746 304292
rect 256602 304240 256608 304292
rect 256660 304280 256666 304292
rect 294598 304280 294604 304292
rect 256660 304252 294604 304280
rect 256660 304240 256666 304252
rect 294598 304240 294604 304252
rect 294656 304240 294662 304292
rect 315850 304240 315856 304292
rect 315908 304280 315914 304292
rect 545114 304280 545120 304292
rect 315908 304252 545120 304280
rect 315908 304240 315914 304252
rect 545114 304240 545120 304252
rect 545172 304240 545178 304292
rect 151722 302880 151728 302932
rect 151780 302920 151786 302932
rect 257062 302920 257068 302932
rect 151780 302892 257068 302920
rect 151780 302880 151786 302892
rect 257062 302880 257068 302892
rect 257120 302880 257126 302932
rect 317138 302880 317144 302932
rect 317196 302920 317202 302932
rect 547138 302920 547144 302932
rect 317196 302892 547144 302920
rect 317196 302880 317202 302892
rect 547138 302880 547144 302892
rect 547196 302880 547202 302932
rect 160002 301452 160008 301504
rect 160060 301492 160066 301504
rect 258074 301492 258080 301504
rect 160060 301464 258080 301492
rect 160060 301452 160066 301464
rect 258074 301452 258080 301464
rect 258132 301452 258138 301504
rect 317230 301452 317236 301504
rect 317288 301492 317294 301504
rect 554774 301492 554780 301504
rect 317288 301464 554780 301492
rect 317288 301452 317294 301464
rect 554774 301452 554780 301464
rect 554832 301452 554838 301504
rect 168282 300092 168288 300144
rect 168340 300132 168346 300144
rect 284938 300132 284944 300144
rect 168340 300104 284944 300132
rect 168340 300092 168346 300104
rect 284938 300092 284944 300104
rect 284996 300092 285002 300144
rect 318610 300092 318616 300144
rect 318668 300132 318674 300144
rect 565078 300132 565084 300144
rect 318668 300104 565084 300132
rect 318668 300092 318674 300104
rect 565078 300092 565084 300104
rect 565136 300092 565142 300144
rect 177942 298732 177948 298784
rect 178000 298772 178006 298784
rect 285766 298772 285772 298784
rect 178000 298744 285772 298772
rect 178000 298732 178006 298744
rect 285766 298732 285772 298744
rect 285824 298732 285830 298784
rect 318702 298732 318708 298784
rect 318760 298772 318766 298784
rect 567838 298772 567844 298784
rect 318760 298744 567844 298772
rect 318760 298732 318766 298744
rect 567838 298732 567844 298744
rect 567896 298732 567902 298784
rect 193122 297372 193128 297424
rect 193180 297412 193186 297424
rect 287790 297412 287796 297424
rect 193180 297384 287796 297412
rect 193180 297372 193186 297384
rect 287790 297372 287796 297384
rect 287848 297372 287854 297424
rect 319898 297372 319904 297424
rect 319956 297412 319962 297424
rect 572714 297412 572720 297424
rect 319956 297384 572720 297412
rect 319956 297372 319962 297384
rect 572714 297372 572720 297384
rect 572772 297372 572778 297424
rect 195882 295944 195888 295996
rect 195940 295984 195946 295996
rect 287698 295984 287704 295996
rect 195940 295956 287704 295984
rect 195940 295944 195946 295956
rect 287698 295944 287704 295956
rect 287756 295944 287762 295996
rect 319990 295944 319996 295996
rect 320048 295984 320054 295996
rect 576118 295984 576124 295996
rect 320048 295956 576124 295984
rect 320048 295944 320054 295956
rect 576118 295944 576124 295956
rect 576176 295944 576182 295996
rect 132402 294584 132408 294636
rect 132460 294624 132466 294636
rect 268378 294624 268384 294636
rect 132460 294596 268384 294624
rect 132460 294584 132466 294596
rect 268378 294584 268384 294596
rect 268436 294584 268442 294636
rect 202782 293224 202788 293276
rect 202840 293264 202846 293276
rect 288618 293264 288624 293276
rect 202840 293236 288624 293264
rect 202840 293224 202846 293236
rect 288618 293224 288624 293236
rect 288676 293224 288682 293276
rect 211062 291796 211068 291848
rect 211120 291836 211126 291848
rect 289998 291836 290004 291848
rect 211120 291808 290004 291836
rect 211120 291796 211126 291808
rect 289998 291796 290004 291808
rect 290056 291796 290062 291848
rect 213822 290436 213828 290488
rect 213880 290476 213886 290488
rect 289906 290476 289912 290488
rect 213880 290448 289912 290476
rect 213880 290436 213886 290448
rect 289906 290436 289912 290448
rect 289964 290436 289970 290488
rect 229002 289144 229008 289196
rect 229060 289184 229066 289196
rect 291930 289184 291936 289196
rect 229060 289156 291936 289184
rect 229060 289144 229066 289156
rect 291930 289144 291936 289156
rect 291988 289144 291994 289196
rect 93762 289076 93768 289128
rect 93820 289116 93826 289128
rect 243078 289116 243084 289128
rect 93820 289088 243084 289116
rect 93820 289076 93826 289088
rect 243078 289076 243084 289088
rect 243136 289076 243142 289128
rect 139302 287648 139308 287700
rect 139360 287688 139366 287700
rect 282086 287688 282092 287700
rect 139360 287660 282092 287688
rect 139360 287648 139366 287660
rect 282086 287648 282092 287660
rect 282144 287648 282150 287700
rect 141970 286288 141976 286340
rect 142028 286328 142034 286340
rect 281718 286328 281724 286340
rect 142028 286300 281724 286328
rect 142028 286288 142034 286300
rect 281718 286288 281724 286300
rect 281776 286288 281782 286340
rect 146202 284928 146208 284980
rect 146260 284968 146266 284980
rect 283098 284968 283104 284980
rect 146260 284940 283104 284968
rect 146260 284928 146266 284940
rect 283098 284928 283104 284940
rect 283156 284928 283162 284980
rect 150342 283568 150348 283620
rect 150400 283608 150406 283620
rect 283006 283608 283012 283620
rect 150400 283580 283012 283608
rect 150400 283568 150406 283580
rect 283006 283568 283012 283580
rect 283064 283568 283070 283620
rect 2038 282140 2044 282192
rect 2096 282180 2102 282192
rect 240318 282180 240324 282192
rect 2096 282152 240324 282180
rect 2096 282140 2102 282152
rect 240318 282140 240324 282152
rect 240376 282140 240382 282192
rect 3418 280780 3424 280832
rect 3476 280820 3482 280832
rect 240502 280820 240508 280832
rect 3476 280792 240508 280820
rect 3476 280780 3482 280792
rect 240502 280780 240508 280792
rect 240560 280780 240566 280832
rect 3142 280100 3148 280152
rect 3200 280140 3206 280152
rect 6178 280140 6184 280152
rect 3200 280112 6184 280140
rect 3200 280100 3206 280112
rect 6178 280100 6184 280112
rect 6236 280100 6242 280152
rect 14458 279420 14464 279472
rect 14516 279460 14522 279472
rect 249978 279460 249984 279472
rect 14516 279432 249984 279460
rect 14516 279420 14522 279432
rect 249978 279420 249984 279432
rect 250036 279420 250042 279472
rect 62022 277992 62028 278044
rect 62080 278032 62086 278044
rect 247218 278032 247224 278044
rect 62080 278004 247224 278032
rect 62080 277992 62086 278004
rect 247218 277992 247224 278004
rect 247276 277992 247282 278044
rect 64782 276632 64788 276684
rect 64840 276672 64846 276684
rect 247678 276672 247684 276684
rect 64840 276644 247684 276672
rect 64840 276632 64846 276644
rect 247678 276632 247684 276644
rect 247736 276632 247742 276684
rect 334618 275952 334624 276004
rect 334676 275992 334682 276004
rect 580166 275992 580172 276004
rect 334676 275964 580172 275992
rect 334676 275952 334682 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 73062 275272 73068 275324
rect 73120 275312 73126 275324
rect 248598 275312 248604 275324
rect 73120 275284 248604 275312
rect 73120 275272 73126 275284
rect 248598 275272 248604 275284
rect 248656 275272 248662 275324
rect 75822 273912 75828 273964
rect 75880 273952 75886 273964
rect 248506 273952 248512 273964
rect 75880 273924 248512 273952
rect 75880 273912 75886 273924
rect 248506 273912 248512 273924
rect 248564 273912 248570 273964
rect 82722 272484 82728 272536
rect 82780 272524 82786 272536
rect 249886 272524 249892 272536
rect 82780 272496 249892 272524
rect 82780 272484 82786 272496
rect 249886 272484 249892 272496
rect 249944 272484 249950 272536
rect 91002 271124 91008 271176
rect 91060 271164 91066 271176
rect 241514 271164 241520 271176
rect 91060 271136 241520 271164
rect 91060 271124 91066 271136
rect 241514 271124 241520 271136
rect 241572 271124 241578 271176
rect 97902 269764 97908 269816
rect 97960 269804 97966 269816
rect 243262 269804 243268 269816
rect 97960 269776 243268 269804
rect 97960 269764 97966 269776
rect 243262 269764 243268 269776
rect 243320 269764 243326 269816
rect 107562 268336 107568 268388
rect 107620 268376 107626 268388
rect 244458 268376 244464 268388
rect 107620 268348 244464 268376
rect 107620 268336 107626 268348
rect 244458 268336 244464 268348
rect 244516 268336 244522 268388
rect 2866 266296 2872 266348
rect 2924 266336 2930 266348
rect 46198 266336 46204 266348
rect 2924 266308 46204 266336
rect 2924 266296 2930 266308
rect 46198 266296 46204 266308
rect 46256 266296 46262 266348
rect 322658 264868 322664 264920
rect 322716 264908 322722 264920
rect 580166 264908 580172 264920
rect 322716 264880 580172 264908
rect 322716 264868 322722 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 326338 252492 326344 252544
rect 326396 252532 326402 252544
rect 579798 252532 579804 252544
rect 326396 252504 579804 252532
rect 326396 252492 326402 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 277210 251812 277216 251864
rect 277268 251852 277274 251864
rect 325694 251852 325700 251864
rect 277268 251824 325700 251852
rect 277268 251812 277274 251824
rect 325694 251812 325700 251824
rect 325752 251812 325758 251864
rect 3510 237328 3516 237380
rect 3568 237368 3574 237380
rect 238386 237368 238392 237380
rect 3568 237340 238392 237368
rect 3568 237328 3574 237340
rect 238386 237328 238392 237340
rect 238444 237328 238450 237380
rect 322566 229032 322572 229084
rect 322624 229072 322630 229084
rect 580166 229072 580172 229084
rect 322624 229044 580172 229072
rect 322624 229032 322630 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 13078 223564 13084 223576
rect 3200 223536 13084 223564
rect 3200 223524 3206 223536
rect 13078 223524 13084 223536
rect 13136 223524 13142 223576
rect 348418 217948 348424 218000
rect 348476 217988 348482 218000
rect 580166 217988 580172 218000
rect 348476 217960 580172 217988
rect 348476 217948 348482 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 280062 217268 280068 217320
rect 280120 217308 280126 217320
rect 347866 217308 347872 217320
rect 280120 217280 347872 217308
rect 280120 217268 280126 217280
rect 347866 217268 347872 217280
rect 347924 217268 347930 217320
rect 2866 194488 2872 194540
rect 2924 194528 2930 194540
rect 28258 194528 28264 194540
rect 2924 194500 28264 194528
rect 2924 194488 2930 194500
rect 28258 194488 28264 194500
rect 28316 194488 28322 194540
rect 333238 182112 333244 182164
rect 333296 182152 333302 182164
rect 580166 182152 580172 182164
rect 333296 182124 580172 182152
rect 333296 182112 333302 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 57238 180792 57244 180804
rect 3292 180764 57244 180792
rect 3292 180752 3298 180764
rect 57238 180752 57244 180764
rect 57296 180752 57302 180804
rect 322474 171028 322480 171080
rect 322532 171068 322538 171080
rect 580166 171068 580172 171080
rect 322532 171040 580172 171068
rect 322532 171028 322538 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 238294 151756 238300 151768
rect 3200 151728 238300 151756
rect 3200 151716 3206 151728
rect 238294 151716 238300 151728
rect 238352 151716 238358 151768
rect 3510 136552 3516 136604
rect 3568 136592 3574 136604
rect 15838 136592 15844 136604
rect 3568 136564 15844 136592
rect 3568 136552 3574 136564
rect 15838 136552 15844 136564
rect 15896 136552 15902 136604
rect 322382 135192 322388 135244
rect 322440 135232 322446 135244
rect 580166 135232 580172 135244
rect 322440 135204 580172 135232
rect 322440 135192 322446 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 317322 133152 317328 133204
rect 317380 133192 317386 133204
rect 552014 133192 552020 133204
rect 317380 133164 552020 133192
rect 317380 133152 317386 133164
rect 552014 133152 552020 133164
rect 552072 133152 552078 133204
rect 341518 124108 341524 124160
rect 341576 124148 341582 124160
rect 580166 124148 580172 124160
rect 341576 124120 580172 124148
rect 341576 124108 341582 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 384298 111732 384304 111784
rect 384356 111772 384362 111784
rect 579798 111772 579804 111784
rect 384356 111744 579804 111772
rect 384356 111732 384362 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 31018 108984 31024 108996
rect 3292 108956 31024 108984
rect 3292 108944 3298 108956
rect 31018 108944 31024 108956
rect 31076 108944 31082 108996
rect 263502 95888 263508 95940
rect 263560 95928 263566 95940
rect 295518 95928 295524 95940
rect 263560 95900 295524 95928
rect 263560 95888 263566 95900
rect 295518 95888 295524 95900
rect 295576 95888 295582 95940
rect 3510 93780 3516 93832
rect 3568 93820 3574 93832
rect 238110 93820 238116 93832
rect 3568 93792 238116 93820
rect 3568 93780 3574 93792
rect 238110 93780 238116 93792
rect 238168 93780 238174 93832
rect 202690 91740 202696 91792
rect 202748 91780 202754 91792
rect 262214 91780 262220 91792
rect 202748 91752 262220 91780
rect 202748 91740 202754 91752
rect 262214 91740 262220 91752
rect 262272 91740 262278 91792
rect 237282 88952 237288 89004
rect 237340 88992 237346 89004
rect 266446 88992 266452 89004
rect 237340 88964 266452 88992
rect 237340 88952 237346 88964
rect 266446 88952 266452 88964
rect 266504 88952 266510 89004
rect 327718 88272 327724 88324
rect 327776 88312 327782 88324
rect 580166 88312 580172 88324
rect 327776 88284 580172 88312
rect 327776 88272 327782 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 322290 77188 322296 77240
rect 322348 77228 322354 77240
rect 580166 77228 580172 77240
rect 322348 77200 580172 77228
rect 322348 77188 322354 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 238202 64852 238208 64864
rect 3384 64824 238208 64852
rect 3384 64812 3390 64824
rect 238202 64812 238208 64824
rect 238260 64812 238266 64864
rect 406378 64812 406384 64864
rect 406436 64852 406442 64864
rect 579798 64852 579804 64864
rect 406436 64824 579804 64852
rect 406436 64812 406442 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 3050 51008 3056 51060
rect 3108 51048 3114 51060
rect 17218 51048 17224 51060
rect 3108 51020 17224 51048
rect 3108 51008 3114 51020
rect 17218 51008 17224 51020
rect 17276 51008 17282 51060
rect 100662 46180 100668 46232
rect 100720 46220 100726 46232
rect 243170 46220 243176 46232
rect 100720 46192 243176 46220
rect 100720 46180 100726 46192
rect 243170 46180 243176 46192
rect 243228 46180 243234 46232
rect 79962 44820 79968 44872
rect 80020 44860 80026 44872
rect 248414 44860 248420 44872
rect 80020 44832 248420 44860
rect 80020 44820 80026 44832
rect 248414 44820 248420 44832
rect 248472 44820 248478 44872
rect 15838 43392 15844 43444
rect 15896 43432 15902 43444
rect 250070 43432 250076 43444
rect 15896 43404 250076 43432
rect 15896 43392 15902 43404
rect 250070 43392 250076 43404
rect 250128 43392 250134 43444
rect 159910 42032 159916 42084
rect 159968 42072 159974 42084
rect 284570 42072 284576 42084
rect 159968 42044 284576 42072
rect 159968 42032 159974 42044
rect 284570 42032 284576 42044
rect 284628 42032 284634 42084
rect 322198 41352 322204 41404
rect 322256 41392 322262 41404
rect 580166 41392 580172 41404
rect 322256 41364 580172 41392
rect 322256 41352 322262 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 68922 40672 68928 40724
rect 68980 40712 68986 40724
rect 247586 40712 247592 40724
rect 68980 40684 247592 40712
rect 68980 40672 68986 40684
rect 247586 40672 247592 40684
rect 247644 40672 247650 40724
rect 235902 39312 235908 39364
rect 235960 39352 235966 39364
rect 292666 39352 292672 39364
rect 235960 39324 292672 39352
rect 235960 39312 235966 39324
rect 292666 39312 292672 39324
rect 292724 39312 292730 39364
rect 153102 37884 153108 37936
rect 153160 37924 153166 37936
rect 282914 37924 282920 37936
rect 153160 37896 282920 37924
rect 153160 37884 153166 37896
rect 282914 37884 282920 37896
rect 282972 37884 282978 37936
rect 238662 36524 238668 36576
rect 238720 36564 238726 36576
rect 292850 36564 292856 36576
rect 238720 36536 292856 36564
rect 238720 36524 238726 36536
rect 292850 36524 292856 36536
rect 292908 36524 292914 36576
rect 224862 35164 224868 35216
rect 224920 35204 224926 35216
rect 291562 35204 291568 35216
rect 224920 35176 291568 35204
rect 224920 35164 224926 35176
rect 291562 35164 291568 35176
rect 291620 35164 291626 35216
rect 220722 33736 220728 33788
rect 220780 33776 220786 33788
rect 291470 33776 291476 33788
rect 220780 33748 291476 33776
rect 220780 33736 220786 33748
rect 291470 33736 291476 33748
rect 291528 33736 291534 33788
rect 206922 32376 206928 32428
rect 206980 32416 206986 32428
rect 289814 32416 289820 32428
rect 206980 32388 289820 32416
rect 206980 32376 206986 32388
rect 289814 32376 289820 32388
rect 289872 32376 289878 32428
rect 217962 31016 217968 31068
rect 218020 31056 218026 31068
rect 290458 31056 290464 31068
rect 218020 31028 290464 31056
rect 218020 31016 218026 31028
rect 290458 31016 290464 31028
rect 290516 31016 290522 31068
rect 340138 30268 340144 30320
rect 340196 30308 340202 30320
rect 580166 30308 580172 30320
rect 340196 30280 580172 30308
rect 340196 30268 340202 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 249702 29656 249708 29708
rect 249760 29696 249766 29708
rect 294322 29696 294328 29708
rect 249760 29668 294328 29696
rect 249760 29656 249766 29668
rect 294322 29656 294328 29668
rect 294380 29656 294386 29708
rect 137922 29588 137928 29640
rect 137980 29628 137986 29640
rect 254578 29628 254584 29640
rect 137980 29600 254584 29628
rect 137980 29588 137986 29600
rect 254578 29588 254584 29600
rect 254636 29588 254642 29640
rect 200022 28228 200028 28280
rect 200080 28268 200086 28280
rect 279510 28268 279516 28280
rect 200080 28240 279516 28268
rect 200080 28228 200086 28240
rect 279510 28228 279516 28240
rect 279568 28228 279574 28280
rect 255222 26936 255228 26988
rect 255280 26976 255286 26988
rect 268286 26976 268292 26988
rect 255280 26948 268292 26976
rect 255280 26936 255286 26948
rect 268286 26936 268292 26948
rect 268344 26936 268350 26988
rect 135162 26868 135168 26920
rect 135220 26908 135226 26920
rect 258810 26908 258816 26920
rect 135220 26880 258816 26908
rect 135220 26868 135226 26880
rect 258810 26868 258816 26880
rect 258868 26868 258874 26920
rect 184842 25508 184848 25560
rect 184900 25548 184906 25560
rect 287146 25548 287152 25560
rect 184900 25520 287152 25548
rect 184900 25508 184906 25520
rect 287146 25508 287152 25520
rect 287204 25508 287210 25560
rect 188982 24080 188988 24132
rect 189040 24120 189046 24132
rect 287422 24120 287428 24132
rect 189040 24092 287428 24120
rect 189040 24080 189046 24092
rect 287422 24080 287428 24092
rect 287480 24080 287486 24132
rect 182082 22720 182088 22772
rect 182140 22760 182146 22772
rect 286318 22760 286324 22772
rect 182140 22732 286324 22760
rect 182140 22720 182146 22732
rect 286318 22720 286324 22732
rect 286376 22720 286382 22772
rect 2866 22040 2872 22092
rect 2924 22080 2930 22092
rect 33778 22080 33784 22092
rect 2924 22052 33784 22080
rect 2924 22040 2930 22052
rect 33778 22040 33784 22052
rect 33836 22040 33842 22092
rect 175182 21360 175188 21412
rect 175240 21400 175246 21412
rect 285858 21400 285864 21412
rect 175240 21372 285864 21400
rect 175240 21360 175246 21372
rect 285858 21360 285864 21372
rect 285916 21360 285922 21412
rect 164142 19932 164148 19984
rect 164200 19972 164206 19984
rect 279418 19972 279424 19984
rect 164200 19944 279424 19972
rect 164200 19932 164206 19944
rect 279418 19932 279424 19944
rect 279476 19932 279482 19984
rect 171042 18572 171048 18624
rect 171100 18612 171106 18624
rect 276658 18612 276664 18624
rect 171100 18584 276664 18612
rect 171100 18572 171106 18584
rect 276658 18572 276664 18584
rect 276716 18572 276722 18624
rect 277302 18572 277308 18624
rect 277360 18612 277366 18624
rect 318794 18612 318800 18624
rect 277360 18584 318800 18612
rect 277360 18572 277366 18584
rect 318794 18572 318800 18584
rect 318852 18572 318858 18624
rect 429838 17892 429844 17944
rect 429896 17932 429902 17944
rect 579798 17932 579804 17944
rect 429896 17904 579804 17932
rect 429896 17892 429902 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 155862 17212 155868 17264
rect 155920 17252 155926 17264
rect 256970 17252 256976 17264
rect 155920 17224 256976 17252
rect 155920 17212 155926 17224
rect 256970 17212 256976 17224
rect 257028 17212 257034 17264
rect 274358 17212 274364 17264
rect 274416 17252 274422 17264
rect 300854 17252 300860 17264
rect 274416 17224 300860 17252
rect 274416 17212 274422 17224
rect 300854 17212 300860 17224
rect 300912 17212 300918 17264
rect 191742 15852 191748 15904
rect 191800 15892 191806 15904
rect 261110 15892 261116 15904
rect 191800 15864 261116 15892
rect 191800 15852 191806 15864
rect 261110 15852 261116 15864
rect 261168 15852 261174 15904
rect 275830 15852 275836 15904
rect 275888 15892 275894 15904
rect 315758 15892 315764 15904
rect 275888 15864 315764 15892
rect 275888 15852 275894 15864
rect 315758 15852 315764 15864
rect 315816 15852 315822 15904
rect 315942 15852 315948 15904
rect 316000 15892 316006 15904
rect 541710 15892 541716 15904
rect 316000 15864 541716 15892
rect 316000 15852 316006 15864
rect 541710 15852 541716 15864
rect 541768 15852 541774 15904
rect 148962 14424 148968 14476
rect 149020 14464 149026 14476
rect 255958 14464 255964 14476
rect 149020 14436 255964 14464
rect 149020 14424 149026 14436
rect 255958 14424 255964 14436
rect 256016 14424 256022 14476
rect 275738 14424 275744 14476
rect 275796 14464 275802 14476
rect 312170 14464 312176 14476
rect 275796 14436 312176 14464
rect 275796 14424 275802 14436
rect 312170 14424 312176 14436
rect 312228 14424 312234 14476
rect 313182 14424 313188 14476
rect 313240 14464 313246 14476
rect 520274 14464 520280 14476
rect 313240 14436 520280 14464
rect 313240 14424 313246 14436
rect 520274 14424 520280 14436
rect 520332 14424 520338 14476
rect 55122 13064 55128 13116
rect 55180 13104 55186 13116
rect 229738 13104 229744 13116
rect 55180 13076 229744 13104
rect 55180 13064 55186 13076
rect 229738 13064 229744 13076
rect 229796 13064 229802 13116
rect 230106 13064 230112 13116
rect 230164 13104 230170 13116
rect 265434 13104 265440 13116
rect 230164 13076 265440 13104
rect 230164 13064 230170 13076
rect 265434 13064 265440 13076
rect 265492 13064 265498 13116
rect 274450 13064 274456 13116
rect 274508 13104 274514 13116
rect 294322 13104 294328 13116
rect 274508 13076 294328 13104
rect 274508 13064 274514 13076
rect 294322 13064 294328 13076
rect 294380 13064 294386 13116
rect 272978 11772 272984 11824
rect 273036 11812 273042 11824
rect 290734 11812 290740 11824
rect 273036 11784 290740 11812
rect 273036 11772 273042 11784
rect 290734 11772 290740 11784
rect 290792 11772 290798 11824
rect 131022 11704 131028 11756
rect 131080 11744 131086 11756
rect 231118 11744 231124 11756
rect 131080 11716 231124 11744
rect 131080 11704 131086 11716
rect 231118 11704 231124 11716
rect 231176 11704 231182 11756
rect 242802 11704 242808 11756
rect 242860 11744 242866 11756
rect 294046 11744 294052 11756
rect 242860 11716 294052 11744
rect 242860 11704 242866 11716
rect 294046 11704 294052 11716
rect 294104 11704 294110 11756
rect 157242 10276 157248 10328
rect 157300 10316 157306 10328
rect 284478 10316 284484 10328
rect 157300 10288 284484 10316
rect 157300 10276 157306 10288
rect 284478 10276 284484 10288
rect 284536 10276 284542 10328
rect 320910 10276 320916 10328
rect 320968 10316 320974 10328
rect 531038 10316 531044 10328
rect 320968 10288 531044 10316
rect 320968 10276 320974 10288
rect 531038 10276 531044 10288
rect 531096 10276 531102 10328
rect 258626 9596 258632 9648
rect 258684 9636 258690 9648
rect 261478 9636 261484 9648
rect 258684 9608 261484 9636
rect 258684 9596 258690 9608
rect 261478 9596 261484 9608
rect 261536 9596 261542 9648
rect 271690 9596 271696 9648
rect 271748 9636 271754 9648
rect 276474 9636 276480 9648
rect 271748 9608 276480 9636
rect 271748 9596 271754 9608
rect 276474 9596 276480 9608
rect 276532 9596 276538 9648
rect 320818 9596 320824 9648
rect 320876 9636 320882 9648
rect 322842 9636 322848 9648
rect 320876 9608 322848 9636
rect 320876 9596 320882 9608
rect 322842 9596 322848 9608
rect 322900 9596 322906 9648
rect 247954 8984 247960 9036
rect 248012 9024 248018 9036
rect 258718 9024 258724 9036
rect 248012 8996 258724 9024
rect 248012 8984 248018 8996
rect 258718 8984 258724 8996
rect 258776 8984 258782 9036
rect 183738 8916 183744 8968
rect 183796 8956 183802 8968
rect 232498 8956 232504 8968
rect 183796 8928 232504 8956
rect 183796 8916 183802 8928
rect 232498 8916 232504 8928
rect 232556 8916 232562 8968
rect 274542 8916 274548 8968
rect 274600 8956 274606 8968
rect 297910 8956 297916 8968
rect 274600 8928 297916 8956
rect 274600 8916 274606 8928
rect 297910 8916 297916 8928
rect 297968 8916 297974 8968
rect 323578 8916 323584 8968
rect 323636 8956 323642 8968
rect 513190 8956 513196 8968
rect 323636 8928 513196 8956
rect 323636 8916 323642 8928
rect 513190 8916 513196 8928
rect 513248 8916 513254 8968
rect 262214 8304 262220 8356
rect 262272 8344 262278 8356
rect 269206 8344 269212 8356
rect 262272 8316 269212 8344
rect 262272 8304 262278 8316
rect 269206 8304 269212 8316
rect 269264 8304 269270 8356
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 238018 8276 238024 8288
rect 3200 8248 238024 8276
rect 3200 8236 3206 8248
rect 238018 8236 238024 8248
rect 238076 8236 238082 8288
rect 244458 7624 244464 7676
rect 244516 7664 244522 7676
rect 265618 7664 265624 7676
rect 244516 7636 265624 7664
rect 244516 7624 244522 7636
rect 265618 7624 265624 7636
rect 265676 7624 265682 7676
rect 273070 7624 273076 7676
rect 273128 7664 273134 7676
rect 287146 7664 287152 7676
rect 273128 7636 287152 7664
rect 273128 7624 273134 7636
rect 287146 7624 287152 7636
rect 287204 7624 287210 7676
rect 252646 7556 252652 7608
rect 252704 7596 252710 7608
rect 291838 7596 291844 7608
rect 252704 7568 291844 7596
rect 252704 7556 252710 7568
rect 291838 7556 291844 7568
rect 291896 7556 291902 7608
rect 310238 7556 310244 7608
rect 310296 7596 310302 7608
rect 495342 7596 495348 7608
rect 310296 7568 495348 7596
rect 310296 7556 310302 7568
rect 495342 7556 495348 7568
rect 495400 7556 495406 7608
rect 265802 6876 265808 6928
rect 265860 6916 265866 6928
rect 269482 6916 269488 6928
rect 265860 6888 269488 6916
rect 265860 6876 265866 6888
rect 269482 6876 269488 6888
rect 269540 6876 269546 6928
rect 251450 6196 251456 6248
rect 251508 6236 251514 6248
rect 267918 6236 267924 6248
rect 251508 6208 267924 6236
rect 251508 6196 251514 6208
rect 267918 6196 267924 6208
rect 267976 6196 267982 6248
rect 281258 6196 281264 6248
rect 281316 6236 281322 6248
rect 354950 6236 354956 6248
rect 281316 6208 354956 6236
rect 281316 6196 281322 6208
rect 354950 6196 354956 6208
rect 355008 6196 355014 6248
rect 172974 6128 172980 6180
rect 173032 6168 173038 6180
rect 233878 6168 233884 6180
rect 173032 6140 233884 6168
rect 173032 6128 173038 6140
rect 233878 6128 233884 6140
rect 233936 6128 233942 6180
rect 262858 6168 262864 6180
rect 238726 6140 262864 6168
rect 233694 6060 233700 6112
rect 233752 6100 233758 6112
rect 238726 6100 238754 6140
rect 262858 6128 262864 6140
rect 262916 6128 262922 6180
rect 281350 6128 281356 6180
rect 281408 6168 281414 6180
rect 358538 6168 358544 6180
rect 281408 6140 358544 6168
rect 281408 6128 281414 6140
rect 358538 6128 358544 6140
rect 358596 6128 358602 6180
rect 233752 6072 238754 6100
rect 233752 6060 233758 6072
rect 240778 4836 240784 4888
rect 240836 4876 240842 4888
rect 266722 4876 266728 4888
rect 240836 4848 266728 4876
rect 240836 4836 240842 4848
rect 266722 4836 266728 4848
rect 266780 4836 266786 4888
rect 273162 4836 273168 4888
rect 273220 4876 273226 4888
rect 280062 4876 280068 4888
rect 273220 4848 280068 4876
rect 273220 4836 273226 4848
rect 280062 4836 280068 4848
rect 280120 4836 280126 4888
rect 165890 4768 165896 4820
rect 165948 4808 165954 4820
rect 236638 4808 236644 4820
rect 165948 4780 236644 4808
rect 165948 4768 165954 4780
rect 236638 4768 236644 4780
rect 236696 4768 236702 4820
rect 245562 4768 245568 4820
rect 245620 4808 245626 4820
rect 293954 4808 293960 4820
rect 245620 4780 293960 4808
rect 245620 4768 245626 4780
rect 293954 4768 293960 4780
rect 294012 4768 294018 4820
rect 308950 4768 308956 4820
rect 309008 4808 309014 4820
rect 484578 4808 484584 4820
rect 309008 4780 484584 4808
rect 309008 4768 309014 4780
rect 484578 4768 484584 4780
rect 484636 4768 484642 4820
rect 271782 4156 271788 4208
rect 271840 4196 271846 4208
rect 272886 4196 272892 4208
rect 271840 4168 272892 4196
rect 271840 4156 271846 4168
rect 272886 4156 272892 4168
rect 272944 4156 272950 4208
rect 280798 4156 280804 4208
rect 280856 4196 280862 4208
rect 283650 4196 283656 4208
rect 280856 4168 283656 4196
rect 280856 4156 280862 4168
rect 283650 4156 283656 4168
rect 283708 4156 283714 4208
rect 312538 4156 312544 4208
rect 312596 4196 312602 4208
rect 313366 4196 313372 4208
rect 312596 4168 313372 4196
rect 312596 4156 312602 4168
rect 313366 4156 313372 4168
rect 313424 4156 313430 4208
rect 127621 4131 127679 4137
rect 127621 4097 127633 4131
rect 127667 4128 127679 4131
rect 245838 4128 245844 4140
rect 127667 4100 245844 4128
rect 127667 4097 127679 4100
rect 127621 4091 127679 4097
rect 245838 4088 245844 4100
rect 245896 4088 245902 4140
rect 311161 4131 311219 4137
rect 311161 4097 311173 4131
rect 311207 4128 311219 4131
rect 324038 4128 324044 4140
rect 311207 4100 324044 4128
rect 311207 4097 311219 4100
rect 311161 4091 311219 4097
rect 324038 4088 324044 4100
rect 324096 4088 324102 4140
rect 547138 4088 547144 4140
rect 547196 4128 547202 4140
rect 548886 4128 548892 4140
rect 547196 4100 548892 4128
rect 547196 4088 547202 4100
rect 548886 4088 548892 4100
rect 548944 4088 548950 4140
rect 576118 4088 576124 4140
rect 576176 4128 576182 4140
rect 577406 4128 577412 4140
rect 576176 4100 577412 4128
rect 576176 4088 576182 4100
rect 577406 4088 577412 4100
rect 577464 4088 577470 4140
rect 114738 4020 114744 4072
rect 114796 4060 114802 4072
rect 244734 4060 244740 4072
rect 114796 4032 244740 4060
rect 114796 4020 114802 4032
rect 244734 4020 244740 4032
rect 244792 4020 244798 4072
rect 295518 4020 295524 4072
rect 295576 4060 295582 4072
rect 299566 4060 299572 4072
rect 295576 4032 299572 4060
rect 295576 4020 295582 4032
rect 299566 4020 299572 4032
rect 299624 4020 299630 4072
rect 304810 4020 304816 4072
rect 304868 4060 304874 4072
rect 327626 4060 327632 4072
rect 304868 4032 327632 4060
rect 304868 4020 304874 4032
rect 327626 4020 327632 4032
rect 327684 4020 327690 4072
rect 111150 3952 111156 4004
rect 111208 3992 111214 4004
rect 244366 3992 244372 4004
rect 111208 3964 244372 3992
rect 111208 3952 111214 3964
rect 244366 3952 244372 3964
rect 244424 3952 244430 4004
rect 248877 3995 248935 4001
rect 248877 3961 248889 3995
rect 248923 3992 248935 3995
rect 252738 3992 252744 4004
rect 248923 3964 252744 3992
rect 248923 3961 248935 3964
rect 248877 3955 248935 3961
rect 252738 3952 252744 3964
rect 252796 3952 252802 4004
rect 291930 3952 291936 4004
rect 291988 3992 291994 4004
rect 299658 3992 299664 4004
rect 291988 3964 299664 3992
rect 291988 3952 291994 3964
rect 299658 3952 299664 3964
rect 299716 3952 299722 4004
rect 304902 3952 304908 4004
rect 304960 3992 304966 4004
rect 331214 3992 331220 4004
rect 304960 3964 331220 3992
rect 304960 3952 304966 3964
rect 331214 3952 331220 3964
rect 331272 3952 331278 4004
rect 46934 3884 46940 3936
rect 46992 3924 46998 3936
rect 253934 3924 253940 3936
rect 46992 3896 253940 3924
rect 46992 3884 46998 3896
rect 253934 3884 253940 3896
rect 253992 3884 253998 3936
rect 288342 3884 288348 3936
rect 288400 3924 288406 3936
rect 299474 3924 299480 3936
rect 288400 3896 299480 3924
rect 288400 3884 288406 3896
rect 299474 3884 299480 3896
rect 299532 3884 299538 3936
rect 303522 3884 303528 3936
rect 303580 3924 303586 3936
rect 311161 3927 311219 3933
rect 311161 3924 311173 3927
rect 303580 3896 311173 3924
rect 303580 3884 303586 3896
rect 311161 3893 311173 3896
rect 311207 3893 311219 3927
rect 311161 3887 311219 3893
rect 311253 3927 311311 3933
rect 311253 3893 311265 3927
rect 311299 3924 311311 3927
rect 334710 3924 334716 3936
rect 311299 3896 334716 3924
rect 311299 3893 311311 3896
rect 311253 3887 311311 3893
rect 334710 3884 334716 3896
rect 334768 3884 334774 3936
rect 43346 3816 43352 3868
rect 43404 3856 43410 3868
rect 252554 3856 252560 3868
rect 43404 3828 252560 3856
rect 43404 3816 43410 3828
rect 252554 3816 252560 3828
rect 252612 3816 252618 3868
rect 284754 3816 284760 3868
rect 284812 3856 284818 3868
rect 298370 3856 298376 3868
rect 284812 3828 298376 3856
rect 284812 3816 284818 3828
rect 298370 3816 298376 3828
rect 298428 3816 298434 3868
rect 306282 3816 306288 3868
rect 306340 3856 306346 3868
rect 338298 3856 338304 3868
rect 306340 3828 338304 3856
rect 306340 3816 306346 3828
rect 338298 3816 338304 3828
rect 338356 3816 338362 3868
rect 39758 3748 39764 3800
rect 39816 3788 39822 3800
rect 252830 3788 252836 3800
rect 39816 3760 252836 3788
rect 39816 3748 39822 3760
rect 252830 3748 252836 3760
rect 252888 3748 252894 3800
rect 281258 3748 281264 3800
rect 281316 3788 281322 3800
rect 298094 3788 298100 3800
rect 281316 3760 298100 3788
rect 281316 3748 281322 3760
rect 298094 3748 298100 3760
rect 298152 3748 298158 3800
rect 306190 3748 306196 3800
rect 306248 3788 306254 3800
rect 341886 3788 341892 3800
rect 306248 3760 341892 3788
rect 306248 3748 306254 3760
rect 341886 3748 341892 3760
rect 341944 3748 341950 3800
rect 36170 3680 36176 3732
rect 36228 3720 36234 3732
rect 248877 3723 248935 3729
rect 248877 3720 248889 3723
rect 36228 3692 248889 3720
rect 36228 3680 36234 3692
rect 248877 3689 248889 3692
rect 248923 3689 248935 3723
rect 248877 3683 248935 3689
rect 248969 3723 249027 3729
rect 248969 3689 248981 3723
rect 249015 3720 249027 3723
rect 251726 3720 251732 3732
rect 249015 3692 251732 3720
rect 249015 3689 249027 3692
rect 248969 3683 249027 3689
rect 251726 3680 251732 3692
rect 251784 3680 251790 3732
rect 277670 3680 277676 3732
rect 277728 3720 277734 3732
rect 298186 3720 298192 3732
rect 277728 3692 298192 3720
rect 277728 3680 277734 3692
rect 298186 3680 298192 3692
rect 298244 3680 298250 3732
rect 304718 3680 304724 3732
rect 304776 3720 304782 3732
rect 311253 3723 311311 3729
rect 311253 3720 311265 3723
rect 304776 3692 311265 3720
rect 304776 3680 304782 3692
rect 311253 3689 311265 3692
rect 311299 3689 311311 3723
rect 311253 3683 311311 3689
rect 311345 3723 311403 3729
rect 311345 3689 311357 3723
rect 311391 3720 311403 3723
rect 349062 3720 349068 3732
rect 311391 3692 349068 3720
rect 311391 3689 311403 3692
rect 311345 3683 311403 3689
rect 349062 3680 349068 3692
rect 349120 3680 349126 3732
rect 32674 3612 32680 3664
rect 32732 3652 32738 3664
rect 251634 3652 251640 3664
rect 32732 3624 251640 3652
rect 32732 3612 32738 3624
rect 251634 3612 251640 3624
rect 251692 3612 251698 3664
rect 281442 3612 281448 3664
rect 281500 3652 281506 3664
rect 363322 3652 363328 3664
rect 281500 3624 363328 3652
rect 281500 3612 281506 3624
rect 363322 3612 363328 3624
rect 363380 3612 363386 3664
rect 29086 3544 29092 3596
rect 29144 3584 29150 3596
rect 248969 3587 249027 3593
rect 248969 3584 248981 3587
rect 29144 3556 248981 3584
rect 29144 3544 29150 3556
rect 248969 3553 248981 3556
rect 249015 3553 249027 3587
rect 251358 3584 251364 3596
rect 248969 3547 249027 3553
rect 249076 3556 251364 3584
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 3418 3516 3424 3528
rect 1728 3488 3424 3516
rect 1728 3476 1734 3488
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 14458 3516 14464 3528
rect 10100 3488 14464 3516
rect 10100 3476 10106 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14826 3476 14832 3528
rect 14884 3516 14890 3528
rect 15838 3516 15844 3528
rect 14884 3488 15844 3516
rect 14884 3476 14890 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 249076 3516 249104 3556
rect 251358 3544 251364 3556
rect 251416 3544 251422 3596
rect 274082 3544 274088 3596
rect 274140 3584 274146 3596
rect 296898 3584 296904 3596
rect 274140 3556 296904 3584
rect 274140 3544 274146 3556
rect 296898 3544 296904 3556
rect 296956 3544 296962 3596
rect 307570 3544 307576 3596
rect 307628 3584 307634 3596
rect 311345 3587 311403 3593
rect 311345 3584 311357 3587
rect 307628 3556 311357 3584
rect 307628 3544 307634 3556
rect 311345 3553 311357 3556
rect 311391 3553 311403 3587
rect 311345 3547 311403 3553
rect 311437 3587 311495 3593
rect 311437 3553 311449 3587
rect 311483 3584 311495 3587
rect 473906 3584 473912 3596
rect 311483 3556 473912 3584
rect 311483 3553 311495 3556
rect 311437 3547 311495 3553
rect 473906 3544 473912 3556
rect 473964 3544 473970 3596
rect 24360 3488 249104 3516
rect 24360 3476 24366 3488
rect 249150 3476 249156 3528
rect 249208 3516 249214 3528
rect 249702 3516 249708 3528
rect 249208 3488 249708 3516
rect 249208 3476 249214 3488
rect 249702 3476 249708 3488
rect 249760 3476 249766 3528
rect 259822 3476 259828 3528
rect 259880 3516 259886 3528
rect 260742 3516 260748 3528
rect 259880 3488 260748 3516
rect 259880 3476 259886 3488
rect 260742 3476 260748 3488
rect 260800 3476 260806 3528
rect 269298 3476 269304 3528
rect 269356 3516 269362 3528
rect 270402 3516 270408 3528
rect 269356 3488 270408 3516
rect 269356 3476 269362 3488
rect 270402 3476 270408 3488
rect 270460 3476 270466 3528
rect 270494 3476 270500 3528
rect 270552 3516 270558 3528
rect 296806 3516 296812 3528
rect 270552 3488 296812 3516
rect 270552 3476 270558 3488
rect 296806 3476 296812 3488
rect 296864 3476 296870 3528
rect 299106 3476 299112 3528
rect 299164 3516 299170 3528
rect 299750 3516 299756 3528
rect 299164 3488 299756 3516
rect 299164 3476 299170 3488
rect 299750 3476 299756 3488
rect 299808 3476 299814 3528
rect 302050 3476 302056 3528
rect 302108 3516 302114 3528
rect 302602 3516 302608 3528
rect 302108 3488 302608 3516
rect 302108 3476 302114 3488
rect 302602 3476 302608 3488
rect 302660 3476 302666 3528
rect 309042 3476 309048 3528
rect 309100 3516 309106 3528
rect 481082 3516 481088 3528
rect 309100 3488 481088 3516
rect 309100 3476 309106 3488
rect 481082 3476 481088 3488
rect 481140 3476 481146 3528
rect 536834 3476 536840 3528
rect 536892 3516 536898 3528
rect 538122 3516 538128 3528
rect 536892 3488 538128 3516
rect 536892 3476 536898 3488
rect 538122 3476 538128 3488
rect 538180 3476 538186 3528
rect 558178 3476 558184 3528
rect 558236 3516 558242 3528
rect 559558 3516 559564 3528
rect 558236 3488 559564 3516
rect 558236 3476 558242 3488
rect 559558 3476 559564 3488
rect 559616 3476 559622 3528
rect 565078 3476 565084 3528
rect 565136 3516 565142 3528
rect 566734 3516 566740 3528
rect 565136 3488 566740 3516
rect 565136 3476 565142 3488
rect 566734 3476 566740 3488
rect 566792 3476 566798 3528
rect 567838 3476 567844 3528
rect 567896 3516 567902 3528
rect 570230 3516 570236 3528
rect 567896 3488 570236 3516
rect 567896 3476 567902 3488
rect 570230 3476 570236 3488
rect 570288 3476 570294 3528
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 10318 3448 10324 3460
rect 2924 3420 10324 3448
rect 2924 3408 2930 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 19518 3408 19524 3460
rect 19576 3448 19582 3460
rect 251266 3448 251272 3460
rect 19576 3420 251272 3448
rect 19576 3408 19582 3420
rect 251266 3408 251272 3420
rect 251324 3408 251330 3460
rect 266998 3408 267004 3460
rect 267056 3448 267062 3460
rect 296714 3448 296720 3460
rect 267056 3420 296720 3448
rect 267056 3408 267062 3420
rect 296714 3408 296720 3420
rect 296772 3408 296778 3460
rect 303430 3408 303436 3460
rect 303488 3448 303494 3460
rect 316954 3448 316960 3460
rect 303488 3420 316960 3448
rect 303488 3408 303494 3420
rect 316954 3408 316960 3420
rect 317012 3408 317018 3460
rect 320082 3408 320088 3460
rect 320140 3448 320146 3460
rect 580994 3448 581000 3460
rect 320140 3420 581000 3448
rect 320140 3408 320146 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 566 3340 572 3392
rect 624 3380 630 3392
rect 2038 3380 2044 3392
rect 624 3352 2044 3380
rect 624 3340 630 3352
rect 2038 3340 2044 3352
rect 2096 3340 2102 3392
rect 50522 3340 50528 3392
rect 50580 3380 50586 3392
rect 50982 3380 50988 3392
rect 50580 3352 50988 3380
rect 50580 3340 50586 3352
rect 50982 3340 50988 3352
rect 51040 3340 51046 3392
rect 54018 3340 54024 3392
rect 54076 3380 54082 3392
rect 55122 3380 55128 3392
rect 54076 3352 55128 3380
rect 54076 3340 54082 3352
rect 55122 3340 55128 3352
rect 55180 3340 55186 3392
rect 61194 3340 61200 3392
rect 61252 3380 61258 3392
rect 62022 3380 62028 3392
rect 61252 3352 62028 3380
rect 61252 3340 61258 3352
rect 62022 3340 62028 3352
rect 62080 3340 62086 3392
rect 68278 3340 68284 3392
rect 68336 3380 68342 3392
rect 68922 3380 68928 3392
rect 68336 3352 68928 3380
rect 68336 3340 68342 3352
rect 68922 3340 68928 3352
rect 68980 3340 68986 3392
rect 71866 3340 71872 3392
rect 71924 3380 71930 3392
rect 73062 3380 73068 3392
rect 71924 3352 73068 3380
rect 71924 3340 71930 3352
rect 73062 3340 73068 3352
rect 73120 3340 73126 3392
rect 79042 3340 79048 3392
rect 79100 3380 79106 3392
rect 79962 3380 79968 3392
rect 79100 3352 79968 3380
rect 79100 3340 79106 3352
rect 79962 3340 79968 3352
rect 80020 3340 80026 3392
rect 89714 3340 89720 3392
rect 89772 3380 89778 3392
rect 91002 3380 91008 3392
rect 89772 3352 91008 3380
rect 89772 3340 89778 3352
rect 91002 3340 91008 3352
rect 91060 3340 91066 3392
rect 93302 3340 93308 3392
rect 93360 3380 93366 3392
rect 93762 3380 93768 3392
rect 93360 3352 93768 3380
rect 93360 3340 93366 3352
rect 93762 3340 93768 3352
rect 93820 3340 93826 3392
rect 96890 3340 96896 3392
rect 96948 3380 96954 3392
rect 97902 3380 97908 3392
rect 96948 3352 97908 3380
rect 96948 3340 96954 3352
rect 97902 3340 97908 3352
rect 97960 3340 97966 3392
rect 103974 3340 103980 3392
rect 104032 3380 104038 3392
rect 104802 3380 104808 3392
rect 104032 3352 104808 3380
rect 104032 3340 104038 3352
rect 104802 3340 104808 3352
rect 104860 3340 104866 3392
rect 118234 3340 118240 3392
rect 118292 3380 118298 3392
rect 127621 3383 127679 3389
rect 127621 3380 127633 3383
rect 118292 3352 127633 3380
rect 118292 3340 118298 3352
rect 127621 3349 127633 3352
rect 127667 3349 127679 3383
rect 127621 3343 127679 3349
rect 130194 3340 130200 3392
rect 130252 3380 130258 3392
rect 131022 3380 131028 3392
rect 130252 3352 131028 3380
rect 130252 3340 130258 3352
rect 131022 3340 131028 3352
rect 131080 3340 131086 3392
rect 240410 3380 240416 3392
rect 131132 3352 240416 3380
rect 121822 3272 121828 3324
rect 121880 3312 121886 3324
rect 122742 3312 122748 3324
rect 121880 3284 122748 3312
rect 121880 3272 121886 3284
rect 122742 3272 122748 3284
rect 122800 3272 122806 3324
rect 125410 3272 125416 3324
rect 125468 3312 125474 3324
rect 131132 3312 131160 3352
rect 240410 3340 240416 3352
rect 240468 3340 240474 3392
rect 241974 3340 241980 3392
rect 242032 3380 242038 3392
rect 242802 3380 242808 3392
rect 242032 3352 242808 3380
rect 242032 3340 242038 3352
rect 242802 3340 242808 3352
rect 242860 3340 242866 3392
rect 303338 3340 303344 3392
rect 303396 3380 303402 3392
rect 320450 3380 320456 3392
rect 303396 3352 320456 3380
rect 303396 3340 303402 3352
rect 320450 3340 320456 3352
rect 320508 3340 320514 3392
rect 339494 3340 339500 3392
rect 339552 3380 339558 3392
rect 340690 3380 340696 3392
rect 339552 3352 340696 3380
rect 339552 3340 339558 3352
rect 340690 3340 340696 3352
rect 340748 3340 340754 3392
rect 125468 3284 131160 3312
rect 125468 3272 125474 3284
rect 131390 3272 131396 3324
rect 131448 3312 131454 3324
rect 132402 3312 132408 3324
rect 131448 3284 132408 3312
rect 131448 3272 131454 3284
rect 132402 3272 132408 3284
rect 132460 3272 132466 3324
rect 137278 3272 137284 3324
rect 137336 3312 137342 3324
rect 137922 3312 137928 3324
rect 137336 3284 137928 3312
rect 137336 3272 137342 3284
rect 137922 3272 137928 3284
rect 137980 3272 137986 3324
rect 138474 3272 138480 3324
rect 138532 3312 138538 3324
rect 139302 3312 139308 3324
rect 138532 3284 139308 3312
rect 138532 3272 138538 3284
rect 139302 3272 139308 3284
rect 139360 3272 139366 3324
rect 140866 3272 140872 3324
rect 140924 3312 140930 3324
rect 142062 3312 142068 3324
rect 140924 3284 142068 3312
rect 140924 3272 140930 3284
rect 142062 3272 142068 3284
rect 142120 3272 142126 3324
rect 145650 3272 145656 3324
rect 145708 3312 145714 3324
rect 146202 3312 146208 3324
rect 145708 3284 146208 3312
rect 145708 3272 145714 3284
rect 146202 3272 146208 3284
rect 146260 3272 146266 3324
rect 148042 3272 148048 3324
rect 148100 3312 148106 3324
rect 148962 3312 148968 3324
rect 148100 3284 148968 3312
rect 148100 3272 148106 3284
rect 148962 3272 148968 3284
rect 149020 3272 149026 3324
rect 149238 3272 149244 3324
rect 149296 3312 149302 3324
rect 150342 3312 150348 3324
rect 149296 3284 150348 3312
rect 149296 3272 149302 3284
rect 150342 3272 150348 3284
rect 150400 3272 150406 3324
rect 155126 3272 155132 3324
rect 155184 3312 155190 3324
rect 155862 3312 155868 3324
rect 155184 3284 155868 3312
rect 155184 3272 155190 3284
rect 155862 3272 155868 3284
rect 155920 3272 155926 3324
rect 156322 3272 156328 3324
rect 156380 3312 156386 3324
rect 157242 3312 157248 3324
rect 156380 3284 157248 3312
rect 156380 3272 156386 3284
rect 157242 3272 157248 3284
rect 157300 3272 157306 3324
rect 158714 3272 158720 3324
rect 158772 3312 158778 3324
rect 160002 3312 160008 3324
rect 158772 3284 160008 3312
rect 158772 3272 158778 3284
rect 160002 3272 160008 3284
rect 160060 3272 160066 3324
rect 162302 3272 162308 3324
rect 162360 3312 162366 3324
rect 162762 3312 162768 3324
rect 162360 3284 162768 3312
rect 162360 3272 162366 3284
rect 162762 3272 162768 3284
rect 162820 3272 162826 3324
rect 163498 3272 163504 3324
rect 163556 3312 163562 3324
rect 164142 3312 164148 3324
rect 163556 3284 164148 3312
rect 163556 3272 163562 3284
rect 164142 3272 164148 3284
rect 164200 3272 164206 3324
rect 167086 3272 167092 3324
rect 167144 3312 167150 3324
rect 168282 3312 168288 3324
rect 167144 3284 168288 3312
rect 167144 3272 167150 3284
rect 168282 3272 168288 3284
rect 168340 3272 168346 3324
rect 170582 3272 170588 3324
rect 170640 3312 170646 3324
rect 171042 3312 171048 3324
rect 170640 3284 171048 3312
rect 170640 3272 170646 3284
rect 171042 3272 171048 3284
rect 171100 3272 171106 3324
rect 174170 3272 174176 3324
rect 174228 3312 174234 3324
rect 175182 3312 175188 3324
rect 174228 3284 175188 3312
rect 174228 3272 174234 3284
rect 175182 3272 175188 3284
rect 175240 3272 175246 3324
rect 180150 3272 180156 3324
rect 180208 3312 180214 3324
rect 180702 3312 180708 3324
rect 180208 3284 180708 3312
rect 180208 3272 180214 3284
rect 180702 3272 180708 3284
rect 180760 3272 180766 3324
rect 181346 3272 181352 3324
rect 181404 3312 181410 3324
rect 182082 3312 182088 3324
rect 181404 3284 182088 3312
rect 181404 3272 181410 3284
rect 182082 3272 182088 3284
rect 182140 3272 182146 3324
rect 190822 3272 190828 3324
rect 190880 3312 190886 3324
rect 191742 3312 191748 3324
rect 190880 3284 191748 3312
rect 190880 3272 190886 3284
rect 191742 3272 191748 3284
rect 191800 3272 191806 3324
rect 192018 3272 192024 3324
rect 192076 3312 192082 3324
rect 193122 3312 193128 3324
rect 192076 3284 193128 3312
rect 192076 3272 192082 3284
rect 193122 3272 193128 3284
rect 193180 3272 193186 3324
rect 197998 3272 198004 3324
rect 198056 3312 198062 3324
rect 198642 3312 198648 3324
rect 198056 3284 198648 3312
rect 198056 3272 198062 3284
rect 198642 3272 198648 3284
rect 198700 3272 198706 3324
rect 199194 3272 199200 3324
rect 199252 3312 199258 3324
rect 200022 3312 200028 3324
rect 199252 3284 200028 3312
rect 199252 3272 199258 3284
rect 200022 3272 200028 3284
rect 200080 3272 200086 3324
rect 201494 3272 201500 3324
rect 201552 3312 201558 3324
rect 202598 3312 202604 3324
rect 201552 3284 202604 3312
rect 201552 3272 201558 3284
rect 202598 3272 202604 3284
rect 202656 3272 202662 3324
rect 205082 3272 205088 3324
rect 205140 3312 205146 3324
rect 205542 3312 205548 3324
rect 205140 3284 205548 3312
rect 205140 3272 205146 3284
rect 205542 3272 205548 3284
rect 205600 3272 205606 3324
rect 206278 3272 206284 3324
rect 206336 3312 206342 3324
rect 206922 3312 206928 3324
rect 206336 3284 206928 3312
rect 206336 3272 206342 3284
rect 206922 3272 206928 3284
rect 206980 3272 206986 3324
rect 208670 3272 208676 3324
rect 208728 3312 208734 3324
rect 209682 3312 209688 3324
rect 208728 3284 209688 3312
rect 208728 3272 208734 3284
rect 209682 3272 209688 3284
rect 209740 3272 209746 3324
rect 209866 3272 209872 3324
rect 209924 3312 209930 3324
rect 211062 3312 211068 3324
rect 209924 3284 211068 3312
rect 209924 3272 209930 3284
rect 211062 3272 211068 3284
rect 211120 3272 211126 3324
rect 215846 3272 215852 3324
rect 215904 3312 215910 3324
rect 216582 3312 216588 3324
rect 215904 3284 216588 3312
rect 215904 3272 215910 3284
rect 216582 3272 216588 3284
rect 216640 3272 216646 3324
rect 217042 3272 217048 3324
rect 217100 3312 217106 3324
rect 217962 3312 217968 3324
rect 217100 3284 217968 3312
rect 217100 3272 217106 3284
rect 217962 3272 217968 3284
rect 218020 3272 218026 3324
rect 222930 3272 222936 3324
rect 222988 3312 222994 3324
rect 223482 3312 223488 3324
rect 222988 3284 223488 3312
rect 222988 3272 222994 3284
rect 223482 3272 223488 3284
rect 223540 3272 223546 3324
rect 224126 3272 224132 3324
rect 224184 3312 224190 3324
rect 224862 3312 224868 3324
rect 224184 3284 224868 3312
rect 224184 3272 224190 3284
rect 224862 3272 224868 3284
rect 224920 3272 224926 3324
rect 226518 3272 226524 3324
rect 226576 3312 226582 3324
rect 227622 3312 227628 3324
rect 226576 3284 227628 3312
rect 226576 3272 226582 3284
rect 227622 3272 227628 3284
rect 227680 3272 227686 3324
rect 227714 3272 227720 3324
rect 227772 3312 227778 3324
rect 229002 3312 229008 3324
rect 227772 3284 229008 3312
rect 227772 3272 227778 3284
rect 229002 3272 229008 3284
rect 229060 3272 229066 3324
rect 231302 3272 231308 3324
rect 231360 3312 231366 3324
rect 231762 3312 231768 3324
rect 231360 3284 231768 3312
rect 231360 3272 231366 3284
rect 231762 3272 231768 3284
rect 231820 3272 231826 3324
rect 234798 3272 234804 3324
rect 234856 3312 234862 3324
rect 235902 3312 235908 3324
rect 234856 3284 235908 3312
rect 234856 3272 234862 3284
rect 235902 3272 235908 3284
rect 235960 3272 235966 3324
rect 307662 3272 307668 3324
rect 307720 3312 307726 3324
rect 311437 3315 311495 3321
rect 311437 3312 311449 3315
rect 307720 3284 311449 3312
rect 307720 3272 307726 3284
rect 311437 3281 311449 3284
rect 311483 3281 311495 3315
rect 311437 3275 311495 3281
rect 188430 3136 188436 3188
rect 188488 3176 188494 3188
rect 188982 3176 188988 3188
rect 188488 3148 188988 3176
rect 188488 3136 188494 3148
rect 188982 3136 188988 3148
rect 189040 3136 189046 3188
rect 302142 3136 302148 3188
rect 302200 3176 302206 3188
rect 306190 3176 306196 3188
rect 302200 3148 306196 3176
rect 302200 3136 302206 3148
rect 306190 3136 306196 3148
rect 306248 3136 306254 3188
rect 86126 2864 86132 2916
rect 86184 2904 86190 2916
rect 86862 2904 86868 2916
rect 86184 2876 86868 2904
rect 86184 2864 86190 2876
rect 86862 2864 86868 2876
rect 86920 2864 86926 2916
rect 554774 2864 554780 2916
rect 554832 2904 554838 2916
rect 555970 2904 555976 2916
rect 554832 2876 555976 2904
rect 554832 2864 554838 2876
rect 555970 2864 555976 2876
rect 556028 2864 556034 2916
<< via1 >>
rect 256608 700408 256660 700460
rect 348792 700408 348844 700460
rect 251088 700340 251140 700392
rect 413652 700340 413704 700392
rect 291108 700272 291160 700324
rect 462320 700272 462372 700324
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 331220 697552 331272 697604
rect 332508 697552 332560 697604
rect 284944 696940 284996 696992
rect 580172 696940 580224 696992
rect 3424 667904 3476 667956
rect 14464 667904 14516 667956
rect 338764 650020 338816 650072
rect 580172 650020 580224 650072
rect 393964 603100 394016 603152
rect 580172 603100 580224 603152
rect 384304 556180 384356 556232
rect 579804 556180 579856 556232
rect 3332 552032 3384 552084
rect 19984 552032 20036 552084
rect 391204 545096 391256 545148
rect 580172 545096 580224 545148
rect 380164 509260 380216 509312
rect 579804 509260 579856 509312
rect 388444 498176 388496 498228
rect 580172 498176 580224 498228
rect 395344 462340 395396 462392
rect 579804 462340 579856 462392
rect 3148 437452 3200 437504
rect 21364 437452 21416 437504
rect 282276 424940 282328 424992
rect 284944 424940 284996 424992
rect 3148 423648 3200 423700
rect 6184 423648 6236 423700
rect 260012 423512 260064 423564
rect 282920 423512 282972 423564
rect 219348 423444 219400 423496
rect 264428 423444 264480 423496
rect 267648 423444 267700 423496
rect 304448 423444 304500 423496
rect 202788 423376 202840 423428
rect 308956 423376 309008 423428
rect 154488 423308 154540 423360
rect 268936 423308 268988 423360
rect 300032 423308 300084 423360
rect 331220 423308 331272 423360
rect 137928 423240 137980 423292
rect 313372 423240 313424 423292
rect 89628 423172 89680 423224
rect 273352 423172 273404 423224
rect 295616 423172 295668 423224
rect 397460 423172 397512 423224
rect 246672 423104 246724 423156
rect 477500 423104 477552 423156
rect 73068 423036 73120 423088
rect 317788 423036 317840 423088
rect 24768 422968 24820 423020
rect 277768 422968 277820 423020
rect 286692 422968 286744 423020
rect 527180 422968 527232 423020
rect 242256 422900 242308 422952
rect 542360 422900 542412 422952
rect 255596 422424 255648 422476
rect 256608 422424 256660 422476
rect 321836 419432 321888 419484
rect 338764 419432 338816 419484
rect 321836 416712 321888 416764
rect 393964 416712 394016 416764
rect 394056 415420 394108 415472
rect 579620 415420 579672 415472
rect 17224 413992 17276 414044
rect 237380 413992 237432 414044
rect 322204 413924 322256 413976
rect 384304 413924 384356 413976
rect 322204 411204 322256 411256
rect 380164 411204 380216 411256
rect 15844 408484 15896 408536
rect 237380 408484 237432 408536
rect 322020 408416 322072 408468
rect 395344 408416 395396 408468
rect 57244 405696 57296 405748
rect 237380 405696 237432 405748
rect 321836 405628 321888 405680
rect 394056 405628 394108 405680
rect 13084 402976 13136 403028
rect 237380 402976 237432 403028
rect 46204 398828 46256 398880
rect 237380 398828 237432 398880
rect 10416 396040 10468 396092
rect 237380 396040 237432 396092
rect 322204 396040 322256 396092
rect 334624 396040 334676 396092
rect 322480 394612 322532 394664
rect 580264 394612 580316 394664
rect 322480 391892 322532 391944
rect 580356 391892 580408 391944
rect 6184 390464 6236 390516
rect 237380 390464 237432 390516
rect 322480 389104 322532 389156
rect 580448 389104 580500 389156
rect 3884 387744 3936 387796
rect 237380 387744 237432 387796
rect 322480 386316 322532 386368
rect 391204 386316 391256 386368
rect 3792 384956 3844 385008
rect 237380 384956 237432 385008
rect 322480 383596 322532 383648
rect 388444 383596 388496 383648
rect 3608 382168 3660 382220
rect 237380 382168 237432 382220
rect 322480 380808 322532 380860
rect 580540 380808 580592 380860
rect 3516 378088 3568 378140
rect 237380 378088 237432 378140
rect 322480 378088 322532 378140
rect 580632 378088 580684 378140
rect 8208 375300 8260 375352
rect 237380 375300 237432 375352
rect 33784 371220 33836 371272
rect 237380 371220 237432 371272
rect 321836 371220 321888 371272
rect 355324 371220 355376 371272
rect 322204 369792 322256 369844
rect 580172 369792 580224 369844
rect 2964 367004 3016 367056
rect 238300 367004 238352 367056
rect 31024 365712 31076 365764
rect 237380 365712 237432 365764
rect 321836 362924 321888 362976
rect 348424 362924 348476 362976
rect 321836 360204 321888 360256
rect 333244 360204 333296 360256
rect 28264 358776 28316 358828
rect 237380 358776 237432 358828
rect 322296 358708 322348 358760
rect 579988 358708 580040 358760
rect 321652 355104 321704 355156
rect 326344 355104 326396 355156
rect 6184 351908 6236 351960
rect 237380 351908 237432 351960
rect 322020 349120 322072 349172
rect 341524 349120 341576 349172
rect 3608 347692 3660 347744
rect 237380 347692 237432 347744
rect 322020 346400 322072 346452
rect 384304 346400 384356 346452
rect 322296 345040 322348 345092
rect 327724 345040 327776 345092
rect 21364 344972 21416 345024
rect 237380 344972 237432 345024
rect 3700 340824 3752 340876
rect 237380 340824 237432 340876
rect 322296 339464 322348 339516
rect 406384 339464 406436 339516
rect 19984 338036 20036 338088
rect 237380 338036 237432 338088
rect 3424 335248 3476 335300
rect 237380 335248 237432 335300
rect 322112 333956 322164 334008
rect 340144 333956 340196 334008
rect 14464 332528 14516 332580
rect 237380 332528 237432 332580
rect 322112 331236 322164 331288
rect 429844 331236 429896 331288
rect 314384 328312 314436 328364
rect 320916 328312 320968 328364
rect 312360 328176 312412 328228
rect 323584 328176 323636 328228
rect 239404 328108 239456 328160
rect 254124 328108 254176 328160
rect 285864 328108 285916 328160
rect 302608 328108 302660 328160
rect 312544 328108 312596 328160
rect 229744 328040 229796 328092
rect 246396 328040 246448 328092
rect 254492 328040 254544 328092
rect 272524 328040 272576 328092
rect 280804 328040 280856 328092
rect 307024 328040 307076 328092
rect 236644 327972 236696 328024
rect 258540 327972 258592 328024
rect 277400 327972 277452 328024
rect 277676 327972 277728 328024
rect 279516 327972 279568 328024
rect 289084 327972 289136 328024
rect 293960 327972 294012 328024
rect 294328 327972 294380 328024
rect 300952 327972 301004 328024
rect 301872 327972 301924 328024
rect 306196 327972 306248 328024
rect 345020 327972 345072 328024
rect 231124 327904 231176 327956
rect 258724 327904 258776 327956
rect 267924 327904 267976 327956
rect 272064 327904 272116 327956
rect 273168 327904 273220 327956
rect 276940 327904 276992 327956
rect 317604 327904 317656 327956
rect 318432 327904 318484 327956
rect 233884 327836 233936 327888
rect 259460 327836 259512 327888
rect 272892 327836 272944 327888
rect 273076 327836 273128 327888
rect 232504 327768 232556 327820
rect 260840 327768 260892 327820
rect 268936 327768 268988 327820
rect 276664 327768 276716 327820
rect 279792 327836 279844 327888
rect 280068 327836 280120 327888
rect 281724 327836 281776 327888
rect 282552 327836 282604 327888
rect 283012 327836 283064 327888
rect 283380 327836 283432 327888
rect 284944 327836 284996 327888
rect 285772 327836 285824 327888
rect 287796 327836 287848 327888
rect 288440 327836 288492 327888
rect 290464 327836 290516 327888
rect 291200 327836 291252 327888
rect 291936 327836 291988 327888
rect 292672 327836 292724 327888
rect 295524 327836 295576 327888
rect 296352 327836 296404 327888
rect 298100 327836 298152 327888
rect 298376 327836 298428 327888
rect 315212 327836 315264 327888
rect 315764 327836 315816 327888
rect 351920 327836 351972 327888
rect 281540 327768 281592 327820
rect 282920 327768 282972 327820
rect 283748 327768 283800 327820
rect 289912 327768 289964 327820
rect 290740 327768 290792 327820
rect 307484 327768 307536 327820
rect 469220 327768 469272 327820
rect 122748 327700 122800 327752
rect 240692 327700 240744 327752
rect 262864 327632 262916 327684
rect 266360 327632 266412 327684
rect 258816 327564 258868 327616
rect 281816 327700 281868 327752
rect 285772 327700 285824 327752
rect 286600 327700 286652 327752
rect 292672 327700 292724 327752
rect 293132 327700 293184 327752
rect 299572 327700 299624 327752
rect 300032 327700 300084 327752
rect 302976 327700 303028 327752
rect 303436 327700 303488 327752
rect 308220 327700 308272 327752
rect 477500 327700 477552 327752
rect 271328 327632 271380 327684
rect 271788 327632 271840 327684
rect 274088 327632 274140 327684
rect 274548 327632 274600 327684
rect 278964 327632 279016 327684
rect 279792 327632 279844 327684
rect 287704 327632 287756 327684
rect 288624 327632 288676 327684
rect 294604 327632 294656 327684
rect 295616 327632 295668 327684
rect 316408 327632 316460 327684
rect 317144 327632 317196 327684
rect 317972 327632 318024 327684
rect 318524 327632 318576 327684
rect 319260 327632 319312 327684
rect 319904 327632 319956 327684
rect 291844 327564 291896 327616
rect 295340 327564 295392 327616
rect 304172 327564 304224 327616
rect 304816 327564 304868 327616
rect 320824 327564 320876 327616
rect 262036 327496 262088 327548
rect 263600 327496 263652 327548
rect 273720 327496 273772 327548
rect 274456 327496 274508 327548
rect 279424 327496 279476 327548
rect 279884 327496 279936 327548
rect 301320 327496 301372 327548
rect 302056 327496 302108 327548
rect 304632 327496 304684 327548
rect 304908 327496 304960 327548
rect 308680 327496 308732 327548
rect 309048 327496 309100 327548
rect 311440 327496 311492 327548
rect 311716 327496 311768 327548
rect 316776 327496 316828 327548
rect 317328 327496 317380 327548
rect 315580 327428 315632 327480
rect 315948 327428 316000 327480
rect 262956 327360 263008 327412
rect 263876 327360 263928 327412
rect 276572 327360 276624 327412
rect 277308 327360 277360 327412
rect 280620 327360 280672 327412
rect 281264 327360 281316 327412
rect 305460 327360 305512 327412
rect 306288 327360 306340 327412
rect 306656 327360 306708 327412
rect 307576 327360 307628 327412
rect 311072 327360 311124 327412
rect 311624 327360 311676 327412
rect 261944 327292 261996 327344
rect 269120 327292 269172 327344
rect 279424 327292 279476 327344
rect 285036 327292 285088 327344
rect 256240 327088 256292 327140
rect 256700 327088 256752 327140
rect 258356 327088 258408 327140
rect 259828 327088 259880 327140
rect 265624 327088 265676 327140
rect 267740 327088 267792 327140
rect 268384 327088 268436 327140
rect 268936 327088 268988 327140
rect 286324 327088 286376 327140
rect 287152 327088 287204 327140
rect 219348 326408 219400 326460
rect 264980 326408 265032 326460
rect 126888 326340 126940 326392
rect 239404 326340 239456 326392
rect 274916 326340 274968 326392
rect 305092 326340 305144 326392
rect 309324 326340 309376 326392
rect 487160 326340 487212 326392
rect 262404 326272 262456 326324
rect 262496 326068 262548 326120
rect 247316 325864 247368 325916
rect 248604 325907 248656 325916
rect 248604 325873 248613 325907
rect 248613 325873 248647 325907
rect 248647 325873 248656 325907
rect 248604 325864 248656 325873
rect 240416 325728 240468 325780
rect 241060 325728 241112 325780
rect 241520 325728 241572 325780
rect 242348 325728 242400 325780
rect 244372 325728 244424 325780
rect 244740 325728 244792 325780
rect 247592 325728 247644 325780
rect 248052 325728 248104 325780
rect 248420 325728 248472 325780
rect 249248 325728 249300 325780
rect 251640 325728 251692 325780
rect 252100 325728 252152 325780
rect 252560 325728 252612 325780
rect 253296 325728 253348 325780
rect 247316 325660 247368 325712
rect 262312 325660 262364 325712
rect 263048 325660 263100 325712
rect 243360 325592 243412 325644
rect 257160 325592 257212 325644
rect 243268 325388 243320 325440
rect 257068 325388 257120 325440
rect 162768 324912 162820 324964
rect 258264 324912 258316 324964
rect 275008 324912 275060 324964
rect 307760 324912 307812 324964
rect 309416 324912 309468 324964
rect 491300 324912 491352 324964
rect 3240 324232 3292 324284
rect 238484 324232 238536 324284
rect 243176 323620 243228 323672
rect 243544 323620 243596 323672
rect 247224 323620 247276 323672
rect 247408 323620 247460 323672
rect 248604 323663 248656 323672
rect 248604 323629 248613 323663
rect 248613 323629 248647 323663
rect 248647 323629 248656 323663
rect 248604 323620 248656 323629
rect 277492 323620 277544 323672
rect 329840 323620 329892 323672
rect 227628 323552 227680 323604
rect 265164 323552 265216 323604
rect 310612 323552 310664 323604
rect 498200 323552 498252 323604
rect 322756 322872 322808 322924
rect 580172 322872 580224 322924
rect 231768 322260 231820 322312
rect 292764 322260 292816 322312
rect 169668 322192 169720 322244
rect 259000 322192 259052 322244
rect 300952 322192 301004 322244
rect 309140 322192 309192 322244
rect 277400 320900 277452 320952
rect 332600 320900 332652 320952
rect 176568 320832 176620 320884
rect 258356 320832 258408 320884
rect 313372 320832 313424 320884
rect 523040 320832 523092 320884
rect 278044 319472 278096 319524
rect 336740 319472 336792 319524
rect 180708 319404 180760 319456
rect 260196 319404 260248 319456
rect 313556 319404 313608 319456
rect 527180 319404 527232 319456
rect 262220 318996 262272 319048
rect 262588 318996 262640 319048
rect 256976 318792 257028 318844
rect 257344 318792 257396 318844
rect 279792 318112 279844 318164
rect 339500 318112 339552 318164
rect 187608 318044 187660 318096
rect 261024 318044 261076 318096
rect 318432 318044 318484 318096
rect 558184 318044 558236 318096
rect 279884 316752 279936 316804
rect 343640 316752 343692 316804
rect 194508 316684 194560 316736
rect 261392 316684 261444 316736
rect 318524 316684 318576 316736
rect 563060 316684 563112 316736
rect 198648 315256 198700 315308
rect 262404 315256 262456 315308
rect 279976 315256 280028 315308
rect 350540 315256 350592 315308
rect 205548 313964 205600 314016
rect 262312 313964 262364 314016
rect 104808 313896 104860 313948
rect 244280 313896 244332 313948
rect 311624 313896 311676 313948
rect 502340 313896 502392 313948
rect 209688 312604 209740 312656
rect 261576 312604 261628 312656
rect 86868 312536 86920 312588
rect 241888 312536 241940 312588
rect 260748 312536 260800 312588
rect 295708 312536 295760 312588
rect 311716 312536 311768 312588
rect 505100 312536 505152 312588
rect 355324 311788 355376 311840
rect 580172 311788 580224 311840
rect 212448 311176 212500 311228
rect 262956 311176 263008 311228
rect 57888 311108 57940 311160
rect 247316 311108 247368 311160
rect 216588 309816 216640 309868
rect 263876 309816 263928 309868
rect 50988 309748 51040 309800
rect 245936 309748 245988 309800
rect 311532 309748 311584 309800
rect 509240 309748 509292 309800
rect 3332 309068 3384 309120
rect 10416 309068 10468 309120
rect 223488 308456 223540 308508
rect 265072 308456 265124 308508
rect 10324 308388 10376 308440
rect 241612 308388 241664 308440
rect 313096 308388 313148 308440
rect 516140 308388 516192 308440
rect 133788 307028 133840 307080
rect 254492 307028 254544 307080
rect 314568 307028 314620 307080
rect 534080 307028 534132 307080
rect 142068 305600 142120 305652
rect 255412 305600 255464 305652
rect 315764 305600 315816 305652
rect 536840 305600 536892 305652
rect 144828 304240 144880 304292
rect 255688 304240 255740 304292
rect 256608 304240 256660 304292
rect 294604 304240 294656 304292
rect 315856 304240 315908 304292
rect 545120 304240 545172 304292
rect 151728 302880 151780 302932
rect 257068 302880 257120 302932
rect 317144 302880 317196 302932
rect 547144 302880 547196 302932
rect 160008 301452 160060 301504
rect 258080 301452 258132 301504
rect 317236 301452 317288 301504
rect 554780 301452 554832 301504
rect 168288 300092 168340 300144
rect 284944 300092 284996 300144
rect 318616 300092 318668 300144
rect 565084 300092 565136 300144
rect 177948 298732 178000 298784
rect 285772 298732 285824 298784
rect 318708 298732 318760 298784
rect 567844 298732 567896 298784
rect 193128 297372 193180 297424
rect 287796 297372 287848 297424
rect 319904 297372 319956 297424
rect 572720 297372 572772 297424
rect 195888 295944 195940 295996
rect 287704 295944 287756 295996
rect 319996 295944 320048 295996
rect 576124 295944 576176 295996
rect 132408 294584 132460 294636
rect 268384 294584 268436 294636
rect 202788 293224 202840 293276
rect 288624 293224 288676 293276
rect 211068 291796 211120 291848
rect 290004 291796 290056 291848
rect 213828 290436 213880 290488
rect 289912 290436 289964 290488
rect 229008 289144 229060 289196
rect 291936 289144 291988 289196
rect 93768 289076 93820 289128
rect 243084 289076 243136 289128
rect 139308 287648 139360 287700
rect 282092 287648 282144 287700
rect 141976 286288 142028 286340
rect 281724 286288 281776 286340
rect 146208 284928 146260 284980
rect 283104 284928 283156 284980
rect 150348 283568 150400 283620
rect 283012 283568 283064 283620
rect 2044 282140 2096 282192
rect 240324 282140 240376 282192
rect 3424 280780 3476 280832
rect 240508 280780 240560 280832
rect 3148 280100 3200 280152
rect 6184 280100 6236 280152
rect 14464 279420 14516 279472
rect 249984 279420 250036 279472
rect 62028 277992 62080 278044
rect 247224 277992 247276 278044
rect 64788 276632 64840 276684
rect 247684 276632 247736 276684
rect 334624 275952 334676 276004
rect 580172 275952 580224 276004
rect 73068 275272 73120 275324
rect 248604 275272 248656 275324
rect 75828 273912 75880 273964
rect 248512 273912 248564 273964
rect 82728 272484 82780 272536
rect 249892 272484 249944 272536
rect 91008 271124 91060 271176
rect 241520 271124 241572 271176
rect 97908 269764 97960 269816
rect 243268 269764 243320 269816
rect 107568 268336 107620 268388
rect 244464 268336 244516 268388
rect 2872 266296 2924 266348
rect 46204 266296 46256 266348
rect 322664 264868 322716 264920
rect 580172 264868 580224 264920
rect 326344 252492 326396 252544
rect 579804 252492 579856 252544
rect 277216 251812 277268 251864
rect 325700 251812 325752 251864
rect 3516 237328 3568 237380
rect 238392 237328 238444 237380
rect 322572 229032 322624 229084
rect 580172 229032 580224 229084
rect 3148 223524 3200 223576
rect 13084 223524 13136 223576
rect 348424 217948 348476 218000
rect 580172 217948 580224 218000
rect 280068 217268 280120 217320
rect 347872 217268 347924 217320
rect 2872 194488 2924 194540
rect 28264 194488 28316 194540
rect 333244 182112 333296 182164
rect 580172 182112 580224 182164
rect 3240 180752 3292 180804
rect 57244 180752 57296 180804
rect 322480 171028 322532 171080
rect 580172 171028 580224 171080
rect 3148 151716 3200 151768
rect 238300 151716 238352 151768
rect 3516 136552 3568 136604
rect 15844 136552 15896 136604
rect 322388 135192 322440 135244
rect 580172 135192 580224 135244
rect 317328 133152 317380 133204
rect 552020 133152 552072 133204
rect 341524 124108 341576 124160
rect 580172 124108 580224 124160
rect 384304 111732 384356 111784
rect 579804 111732 579856 111784
rect 3240 108944 3292 108996
rect 31024 108944 31076 108996
rect 263508 95888 263560 95940
rect 295524 95888 295576 95940
rect 3516 93780 3568 93832
rect 238116 93780 238168 93832
rect 202696 91740 202748 91792
rect 262220 91740 262272 91792
rect 237288 88952 237340 89004
rect 266452 88952 266504 89004
rect 327724 88272 327776 88324
rect 580172 88272 580224 88324
rect 322296 77188 322348 77240
rect 580172 77188 580224 77240
rect 3332 64812 3384 64864
rect 238208 64812 238260 64864
rect 406384 64812 406436 64864
rect 579804 64812 579856 64864
rect 3056 51008 3108 51060
rect 17224 51008 17276 51060
rect 100668 46180 100720 46232
rect 243176 46180 243228 46232
rect 79968 44820 80020 44872
rect 248420 44820 248472 44872
rect 15844 43392 15896 43444
rect 250076 43392 250128 43444
rect 159916 42032 159968 42084
rect 284576 42032 284628 42084
rect 322204 41352 322256 41404
rect 580172 41352 580224 41404
rect 68928 40672 68980 40724
rect 247592 40672 247644 40724
rect 235908 39312 235960 39364
rect 292672 39312 292724 39364
rect 153108 37884 153160 37936
rect 282920 37884 282972 37936
rect 238668 36524 238720 36576
rect 292856 36524 292908 36576
rect 224868 35164 224920 35216
rect 291568 35164 291620 35216
rect 220728 33736 220780 33788
rect 291476 33736 291528 33788
rect 206928 32376 206980 32428
rect 289820 32376 289872 32428
rect 217968 31016 218020 31068
rect 290464 31016 290516 31068
rect 340144 30268 340196 30320
rect 580172 30268 580224 30320
rect 249708 29656 249760 29708
rect 294328 29656 294380 29708
rect 137928 29588 137980 29640
rect 254584 29588 254636 29640
rect 200028 28228 200080 28280
rect 279516 28228 279568 28280
rect 255228 26936 255280 26988
rect 268292 26936 268344 26988
rect 135168 26868 135220 26920
rect 258816 26868 258868 26920
rect 184848 25508 184900 25560
rect 287152 25508 287204 25560
rect 188988 24080 189040 24132
rect 287428 24080 287480 24132
rect 182088 22720 182140 22772
rect 286324 22720 286376 22772
rect 2872 22040 2924 22092
rect 33784 22040 33836 22092
rect 175188 21360 175240 21412
rect 285864 21360 285916 21412
rect 164148 19932 164200 19984
rect 279424 19932 279476 19984
rect 171048 18572 171100 18624
rect 276664 18572 276716 18624
rect 277308 18572 277360 18624
rect 318800 18572 318852 18624
rect 429844 17892 429896 17944
rect 579804 17892 579856 17944
rect 155868 17212 155920 17264
rect 256976 17212 257028 17264
rect 274364 17212 274416 17264
rect 300860 17212 300912 17264
rect 191748 15852 191800 15904
rect 261116 15852 261168 15904
rect 275836 15852 275888 15904
rect 315764 15852 315816 15904
rect 315948 15852 316000 15904
rect 541716 15852 541768 15904
rect 148968 14424 149020 14476
rect 255964 14424 256016 14476
rect 275744 14424 275796 14476
rect 312176 14424 312228 14476
rect 313188 14424 313240 14476
rect 520280 14424 520332 14476
rect 55128 13064 55180 13116
rect 229744 13064 229796 13116
rect 230112 13064 230164 13116
rect 265440 13064 265492 13116
rect 274456 13064 274508 13116
rect 294328 13064 294380 13116
rect 272984 11772 273036 11824
rect 290740 11772 290792 11824
rect 131028 11704 131080 11756
rect 231124 11704 231176 11756
rect 242808 11704 242860 11756
rect 294052 11704 294104 11756
rect 157248 10276 157300 10328
rect 284484 10276 284536 10328
rect 320916 10276 320968 10328
rect 531044 10276 531096 10328
rect 258632 9596 258684 9648
rect 261484 9596 261536 9648
rect 271696 9596 271748 9648
rect 276480 9596 276532 9648
rect 320824 9596 320876 9648
rect 322848 9596 322900 9648
rect 247960 8984 248012 9036
rect 258724 8984 258776 9036
rect 183744 8916 183796 8968
rect 232504 8916 232556 8968
rect 274548 8916 274600 8968
rect 297916 8916 297968 8968
rect 323584 8916 323636 8968
rect 513196 8916 513248 8968
rect 262220 8304 262272 8356
rect 269212 8304 269264 8356
rect 3148 8236 3200 8288
rect 238024 8236 238076 8288
rect 244464 7624 244516 7676
rect 265624 7624 265676 7676
rect 273076 7624 273128 7676
rect 287152 7624 287204 7676
rect 252652 7556 252704 7608
rect 291844 7556 291896 7608
rect 310244 7556 310296 7608
rect 495348 7556 495400 7608
rect 265808 6876 265860 6928
rect 269488 6876 269540 6928
rect 251456 6196 251508 6248
rect 267924 6196 267976 6248
rect 281264 6196 281316 6248
rect 354956 6196 355008 6248
rect 172980 6128 173032 6180
rect 233884 6128 233936 6180
rect 233700 6060 233752 6112
rect 262864 6128 262916 6180
rect 281356 6128 281408 6180
rect 358544 6128 358596 6180
rect 240784 4836 240836 4888
rect 266728 4836 266780 4888
rect 273168 4836 273220 4888
rect 280068 4836 280120 4888
rect 165896 4768 165948 4820
rect 236644 4768 236696 4820
rect 245568 4768 245620 4820
rect 293960 4768 294012 4820
rect 308956 4768 309008 4820
rect 484584 4768 484636 4820
rect 271788 4156 271840 4208
rect 272892 4156 272944 4208
rect 280804 4156 280856 4208
rect 283656 4156 283708 4208
rect 312544 4156 312596 4208
rect 313372 4156 313424 4208
rect 245844 4088 245896 4140
rect 324044 4088 324096 4140
rect 547144 4088 547196 4140
rect 548892 4088 548944 4140
rect 576124 4088 576176 4140
rect 577412 4088 577464 4140
rect 114744 4020 114796 4072
rect 244740 4020 244792 4072
rect 295524 4020 295576 4072
rect 299572 4020 299624 4072
rect 304816 4020 304868 4072
rect 327632 4020 327684 4072
rect 111156 3952 111208 4004
rect 244372 3952 244424 4004
rect 252744 3952 252796 4004
rect 291936 3952 291988 4004
rect 299664 3952 299716 4004
rect 304908 3952 304960 4004
rect 331220 3952 331272 4004
rect 46940 3884 46992 3936
rect 253940 3884 253992 3936
rect 288348 3884 288400 3936
rect 299480 3884 299532 3936
rect 303528 3884 303580 3936
rect 334716 3884 334768 3936
rect 43352 3816 43404 3868
rect 252560 3816 252612 3868
rect 284760 3816 284812 3868
rect 298376 3816 298428 3868
rect 306288 3816 306340 3868
rect 338304 3816 338356 3868
rect 39764 3748 39816 3800
rect 252836 3748 252888 3800
rect 281264 3748 281316 3800
rect 298100 3748 298152 3800
rect 306196 3748 306248 3800
rect 341892 3748 341944 3800
rect 36176 3680 36228 3732
rect 251732 3680 251784 3732
rect 277676 3680 277728 3732
rect 298192 3680 298244 3732
rect 304724 3680 304776 3732
rect 349068 3680 349120 3732
rect 32680 3612 32732 3664
rect 251640 3612 251692 3664
rect 281448 3612 281500 3664
rect 363328 3612 363380 3664
rect 29092 3544 29144 3596
rect 1676 3476 1728 3528
rect 3424 3476 3476 3528
rect 10048 3476 10100 3528
rect 14464 3476 14516 3528
rect 14832 3476 14884 3528
rect 15844 3476 15896 3528
rect 24308 3476 24360 3528
rect 251364 3544 251416 3596
rect 274088 3544 274140 3596
rect 296904 3544 296956 3596
rect 307576 3544 307628 3596
rect 473912 3544 473964 3596
rect 249156 3476 249208 3528
rect 249708 3476 249760 3528
rect 259828 3476 259880 3528
rect 260748 3476 260800 3528
rect 269304 3476 269356 3528
rect 270408 3476 270460 3528
rect 270500 3476 270552 3528
rect 296812 3476 296864 3528
rect 299112 3476 299164 3528
rect 299756 3476 299808 3528
rect 302056 3476 302108 3528
rect 302608 3476 302660 3528
rect 309048 3476 309100 3528
rect 481088 3476 481140 3528
rect 536840 3476 536892 3528
rect 538128 3476 538180 3528
rect 558184 3476 558236 3528
rect 559564 3476 559616 3528
rect 565084 3476 565136 3528
rect 566740 3476 566792 3528
rect 567844 3476 567896 3528
rect 570236 3476 570288 3528
rect 2872 3408 2924 3460
rect 10324 3408 10376 3460
rect 19524 3408 19576 3460
rect 251272 3408 251324 3460
rect 267004 3408 267056 3460
rect 296720 3408 296772 3460
rect 303436 3408 303488 3460
rect 316960 3408 317012 3460
rect 320088 3408 320140 3460
rect 581000 3408 581052 3460
rect 572 3340 624 3392
rect 2044 3340 2096 3392
rect 50528 3340 50580 3392
rect 50988 3340 51040 3392
rect 54024 3340 54076 3392
rect 55128 3340 55180 3392
rect 61200 3340 61252 3392
rect 62028 3340 62080 3392
rect 68284 3340 68336 3392
rect 68928 3340 68980 3392
rect 71872 3340 71924 3392
rect 73068 3340 73120 3392
rect 79048 3340 79100 3392
rect 79968 3340 80020 3392
rect 89720 3340 89772 3392
rect 91008 3340 91060 3392
rect 93308 3340 93360 3392
rect 93768 3340 93820 3392
rect 96896 3340 96948 3392
rect 97908 3340 97960 3392
rect 103980 3340 104032 3392
rect 104808 3340 104860 3392
rect 118240 3340 118292 3392
rect 130200 3340 130252 3392
rect 131028 3340 131080 3392
rect 121828 3272 121880 3324
rect 122748 3272 122800 3324
rect 125416 3272 125468 3324
rect 240416 3340 240468 3392
rect 241980 3340 242032 3392
rect 242808 3340 242860 3392
rect 303344 3340 303396 3392
rect 320456 3340 320508 3392
rect 339500 3340 339552 3392
rect 340696 3340 340748 3392
rect 131396 3272 131448 3324
rect 132408 3272 132460 3324
rect 137284 3272 137336 3324
rect 137928 3272 137980 3324
rect 138480 3272 138532 3324
rect 139308 3272 139360 3324
rect 140872 3272 140924 3324
rect 142068 3272 142120 3324
rect 145656 3272 145708 3324
rect 146208 3272 146260 3324
rect 148048 3272 148100 3324
rect 148968 3272 149020 3324
rect 149244 3272 149296 3324
rect 150348 3272 150400 3324
rect 155132 3272 155184 3324
rect 155868 3272 155920 3324
rect 156328 3272 156380 3324
rect 157248 3272 157300 3324
rect 158720 3272 158772 3324
rect 160008 3272 160060 3324
rect 162308 3272 162360 3324
rect 162768 3272 162820 3324
rect 163504 3272 163556 3324
rect 164148 3272 164200 3324
rect 167092 3272 167144 3324
rect 168288 3272 168340 3324
rect 170588 3272 170640 3324
rect 171048 3272 171100 3324
rect 174176 3272 174228 3324
rect 175188 3272 175240 3324
rect 180156 3272 180208 3324
rect 180708 3272 180760 3324
rect 181352 3272 181404 3324
rect 182088 3272 182140 3324
rect 190828 3272 190880 3324
rect 191748 3272 191800 3324
rect 192024 3272 192076 3324
rect 193128 3272 193180 3324
rect 198004 3272 198056 3324
rect 198648 3272 198700 3324
rect 199200 3272 199252 3324
rect 200028 3272 200080 3324
rect 201500 3272 201552 3324
rect 202604 3272 202656 3324
rect 205088 3272 205140 3324
rect 205548 3272 205600 3324
rect 206284 3272 206336 3324
rect 206928 3272 206980 3324
rect 208676 3272 208728 3324
rect 209688 3272 209740 3324
rect 209872 3272 209924 3324
rect 211068 3272 211120 3324
rect 215852 3272 215904 3324
rect 216588 3272 216640 3324
rect 217048 3272 217100 3324
rect 217968 3272 218020 3324
rect 222936 3272 222988 3324
rect 223488 3272 223540 3324
rect 224132 3272 224184 3324
rect 224868 3272 224920 3324
rect 226524 3272 226576 3324
rect 227628 3272 227680 3324
rect 227720 3272 227772 3324
rect 229008 3272 229060 3324
rect 231308 3272 231360 3324
rect 231768 3272 231820 3324
rect 234804 3272 234856 3324
rect 235908 3272 235960 3324
rect 307668 3272 307720 3324
rect 188436 3136 188488 3188
rect 188988 3136 189040 3188
rect 302148 3136 302200 3188
rect 306196 3136 306248 3188
rect 86132 2864 86184 2916
rect 86868 2864 86920 2916
rect 554780 2864 554832 2916
rect 555976 2864 556028 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3514 653576 3570 653585
rect 3514 653511 3570 653520
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3330 553072 3386 553081
rect 3330 553007 3386 553016
rect 3344 552090 3372 553007
rect 3332 552084 3384 552090
rect 3332 552026 3384 552032
rect 3146 438016 3202 438025
rect 3146 437951 3202 437960
rect 3160 437510 3188 437951
rect 3148 437504 3200 437510
rect 3148 437446 3200 437452
rect 3146 423736 3202 423745
rect 3146 423671 3148 423680
rect 3200 423671 3202 423680
rect 3148 423642 3200 423648
rect 2964 367056 3016 367062
rect 2964 366998 3016 367004
rect 2976 366217 3004 366998
rect 2962 366208 3018 366217
rect 2962 366143 3018 366152
rect 3436 335306 3464 610399
rect 3528 378146 3556 653511
rect 3606 596048 3662 596057
rect 3606 595983 3662 595992
rect 3620 382226 3648 595983
rect 3790 538656 3846 538665
rect 3790 538591 3846 538600
rect 3698 495544 3754 495553
rect 3698 495479 3754 495488
rect 3608 382220 3660 382226
rect 3608 382162 3660 382168
rect 3606 380624 3662 380633
rect 3606 380559 3662 380568
rect 3516 378140 3568 378146
rect 3516 378082 3568 378088
rect 3620 347750 3648 380559
rect 3608 347744 3660 347750
rect 3608 347686 3660 347692
rect 3712 340882 3740 495479
rect 3804 385014 3832 538591
rect 3882 481128 3938 481137
rect 3882 481063 3938 481072
rect 3896 387802 3924 481063
rect 6184 423700 6236 423706
rect 6184 423642 6236 423648
rect 6196 390522 6224 423642
rect 6184 390516 6236 390522
rect 6184 390458 6236 390464
rect 3884 387796 3936 387802
rect 3884 387738 3936 387744
rect 3792 385008 3844 385014
rect 3792 384950 3844 384956
rect 8220 375358 8248 702406
rect 24320 699718 24348 703520
rect 72988 702434 73016 703520
rect 72988 702406 73108 702434
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 14464 667956 14516 667962
rect 14464 667898 14516 667904
rect 13084 403028 13136 403034
rect 13084 402970 13136 402976
rect 10416 396092 10468 396098
rect 10416 396034 10468 396040
rect 8208 375352 8260 375358
rect 8208 375294 8260 375300
rect 6184 351960 6236 351966
rect 6184 351902 6236 351908
rect 3700 340876 3752 340882
rect 3700 340818 3752 340824
rect 3424 335300 3476 335306
rect 3424 335242 3476 335248
rect 3240 324284 3292 324290
rect 3240 324226 3292 324232
rect 3252 323105 3280 324226
rect 3238 323096 3294 323105
rect 3238 323031 3294 323040
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 2044 282192 2096 282198
rect 2044 282134 2096 282140
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3392 624 3398
rect 572 3334 624 3340
rect 584 480 612 3334
rect 1688 480 1716 3470
rect 2056 3398 2084 282134
rect 3424 280832 3476 280838
rect 3424 280774 3476 280780
rect 3148 280152 3200 280158
rect 3146 280120 3148 280129
rect 3200 280120 3202 280129
rect 3146 280055 3202 280064
rect 2872 266348 2924 266354
rect 2872 266290 2924 266296
rect 2884 265713 2912 266290
rect 2870 265704 2926 265713
rect 2870 265639 2926 265648
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 2872 194540 2924 194546
rect 2872 194482 2924 194488
rect 2884 193905 2912 194482
rect 2870 193896 2926 193905
rect 2870 193831 2926 193840
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3056 51060 3108 51066
rect 3056 51002 3108 51008
rect 3068 50153 3096 51002
rect 3054 50144 3110 50153
rect 3054 50079 3110 50088
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2884 21457 2912 22034
rect 2870 21448 2926 21457
rect 2870 21383 2926 21392
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3160 7177 3188 8230
rect 3146 7168 3202 7177
rect 3146 7103 3202 7112
rect 3436 3534 3464 280774
rect 6196 280158 6224 351902
rect 10428 309126 10456 396034
rect 10416 309120 10468 309126
rect 10416 309062 10468 309068
rect 10324 308440 10376 308446
rect 10324 308382 10376 308388
rect 6184 280152 6236 280158
rect 6184 280094 6236 280100
rect 3516 237380 3568 237386
rect 3516 237322 3568 237328
rect 3528 237017 3556 237322
rect 3514 237008 3570 237017
rect 3514 236943 3570 236952
rect 3516 136604 3568 136610
rect 3516 136546 3568 136552
rect 3528 136377 3556 136546
rect 3514 136368 3570 136377
rect 3514 136303 3570 136312
rect 3516 93832 3568 93838
rect 3516 93774 3568 93780
rect 3528 93265 3556 93774
rect 3514 93256 3570 93265
rect 3514 93191 3570 93200
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2884 480 2912 3402
rect 10060 480 10088 3470
rect 10336 3466 10364 308382
rect 13096 223582 13124 402970
rect 14476 332586 14504 667898
rect 19984 552084 20036 552090
rect 19984 552026 20036 552032
rect 17224 414044 17276 414050
rect 17224 413986 17276 413992
rect 15844 408536 15896 408542
rect 15844 408478 15896 408484
rect 14464 332580 14516 332586
rect 14464 332522 14516 332528
rect 14464 279472 14516 279478
rect 14464 279414 14516 279420
rect 13084 223576 13136 223582
rect 13084 223518 13136 223524
rect 14476 3534 14504 279414
rect 15856 136610 15884 408478
rect 15844 136604 15896 136610
rect 15844 136546 15896 136552
rect 17236 51066 17264 413986
rect 19996 338094 20024 552026
rect 21364 437504 21416 437510
rect 21364 437446 21416 437452
rect 21376 345030 21404 437446
rect 24780 423026 24808 699654
rect 73080 423094 73108 702406
rect 89180 699718 89208 703520
rect 137848 702434 137876 703520
rect 154132 702434 154160 703520
rect 137848 702406 137968 702434
rect 154132 702406 154528 702434
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 89640 423230 89668 699654
rect 137940 423298 137968 702406
rect 154500 423366 154528 702406
rect 202800 423434 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 219360 423502 219388 702406
rect 256608 700460 256660 700466
rect 256608 700402 256660 700408
rect 251088 700392 251140 700398
rect 251088 700334 251140 700340
rect 219348 423496 219400 423502
rect 219348 423438 219400 423444
rect 202788 423428 202840 423434
rect 202788 423370 202840 423376
rect 154488 423360 154540 423366
rect 154488 423302 154540 423308
rect 137928 423292 137980 423298
rect 137928 423234 137980 423240
rect 89628 423224 89680 423230
rect 89628 423166 89680 423172
rect 246672 423156 246724 423162
rect 246672 423098 246724 423104
rect 73068 423088 73120 423094
rect 73068 423030 73120 423036
rect 24768 423020 24820 423026
rect 24768 422962 24820 422968
rect 242256 422952 242308 422958
rect 242256 422894 242308 422900
rect 242268 419900 242296 422894
rect 246684 419900 246712 423098
rect 251100 419900 251128 700334
rect 256620 422482 256648 700402
rect 260012 423564 260064 423570
rect 260012 423506 260064 423512
rect 255596 422476 255648 422482
rect 255596 422418 255648 422424
rect 256608 422476 256660 422482
rect 256608 422418 256660 422424
rect 255608 419900 255636 422418
rect 260024 419900 260052 423506
rect 267660 423502 267688 703520
rect 283852 683114 283880 703520
rect 291108 700324 291160 700330
rect 291108 700266 291160 700272
rect 284944 696992 284996 696998
rect 284944 696934 284996 696940
rect 282932 683086 283880 683114
rect 282276 424992 282328 424998
rect 282276 424934 282328 424940
rect 264428 423496 264480 423502
rect 264428 423438 264480 423444
rect 267648 423496 267700 423502
rect 267648 423438 267700 423444
rect 264440 419900 264468 423438
rect 268936 423360 268988 423366
rect 268936 423302 268988 423308
rect 268948 419900 268976 423302
rect 273352 423224 273404 423230
rect 273352 423166 273404 423172
rect 273364 419900 273392 423166
rect 277768 423020 277820 423026
rect 277768 422962 277820 422968
rect 277780 419900 277808 422962
rect 282288 419900 282316 424934
rect 282932 423570 282960 683086
rect 284956 424998 284984 696934
rect 284944 424992 284996 424998
rect 284944 424934 284996 424940
rect 282920 423564 282972 423570
rect 282920 423506 282972 423512
rect 286692 423020 286744 423026
rect 286692 422962 286744 422968
rect 286704 419900 286732 422962
rect 291120 419900 291148 700266
rect 332520 697610 332548 703520
rect 348804 700466 348832 703520
rect 348792 700460 348844 700466
rect 348792 700402 348844 700408
rect 331220 697604 331272 697610
rect 331220 697546 331272 697552
rect 332508 697604 332560 697610
rect 332508 697546 332560 697552
rect 304448 423496 304500 423502
rect 304448 423438 304500 423444
rect 300032 423360 300084 423366
rect 300032 423302 300084 423308
rect 295616 423224 295668 423230
rect 295616 423166 295668 423172
rect 295628 419900 295656 423166
rect 300044 419900 300072 423302
rect 304460 419900 304488 423438
rect 308956 423428 309008 423434
rect 308956 423370 309008 423376
rect 308968 419900 308996 423370
rect 331232 423366 331260 697546
rect 338764 650072 338816 650078
rect 338764 650014 338816 650020
rect 331220 423360 331272 423366
rect 331220 423302 331272 423308
rect 313372 423292 313424 423298
rect 313372 423234 313424 423240
rect 313384 419900 313412 423234
rect 317788 423088 317840 423094
rect 317788 423030 317840 423036
rect 317800 419900 317828 423030
rect 338776 419490 338804 650014
rect 393964 603152 394016 603158
rect 393964 603094 394016 603100
rect 384304 556232 384356 556238
rect 384304 556174 384356 556180
rect 380164 509312 380216 509318
rect 380164 509254 380216 509260
rect 321836 419484 321888 419490
rect 321836 419426 321888 419432
rect 338764 419484 338816 419490
rect 338764 419426 338816 419432
rect 321848 419121 321876 419426
rect 321834 419112 321890 419121
rect 321834 419047 321890 419056
rect 238022 418296 238078 418305
rect 238022 418231 238078 418240
rect 237378 414760 237434 414769
rect 237378 414695 237434 414704
rect 237392 414050 237420 414695
rect 237380 414044 237432 414050
rect 237380 413986 237432 413992
rect 237378 408776 237434 408785
rect 237378 408711 237434 408720
rect 237392 408542 237420 408711
rect 237380 408536 237432 408542
rect 237380 408478 237432 408484
rect 237378 405784 237434 405793
rect 57244 405748 57296 405754
rect 237378 405719 237380 405728
rect 57244 405690 57296 405696
rect 237432 405719 237434 405728
rect 237380 405690 237432 405696
rect 46204 398880 46256 398886
rect 46204 398822 46256 398828
rect 33784 371272 33836 371278
rect 33784 371214 33836 371220
rect 31024 365764 31076 365770
rect 31024 365706 31076 365712
rect 28264 358828 28316 358834
rect 28264 358770 28316 358776
rect 21364 345024 21416 345030
rect 21364 344966 21416 344972
rect 19984 338088 20036 338094
rect 19984 338030 20036 338036
rect 28276 194546 28304 358770
rect 28264 194540 28316 194546
rect 28264 194482 28316 194488
rect 31036 109002 31064 365706
rect 31024 108996 31076 109002
rect 31024 108938 31076 108944
rect 17224 51060 17276 51066
rect 17224 51002 17276 51008
rect 15844 43444 15896 43450
rect 15844 43386 15896 43392
rect 15856 3534 15884 43386
rect 33796 22098 33824 371214
rect 46216 266354 46244 398822
rect 50988 309800 51040 309806
rect 50988 309742 51040 309748
rect 46204 266348 46256 266354
rect 46204 266290 46256 266296
rect 33784 22092 33836 22098
rect 33784 22034 33836 22040
rect 46940 3936 46992 3942
rect 46940 3878 46992 3884
rect 43352 3868 43404 3874
rect 43352 3810 43404 3816
rect 39764 3800 39816 3806
rect 39764 3742 39816 3748
rect 36176 3732 36228 3738
rect 36176 3674 36228 3680
rect 32680 3664 32732 3670
rect 32680 3606 32732 3612
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 14844 480 14872 3470
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19536 480 19564 3402
rect 24320 480 24348 3470
rect 29104 480 29132 3538
rect 32692 480 32720 3606
rect 36188 480 36216 3674
rect 39776 480 39804 3742
rect 43364 480 43392 3810
rect 46952 480 46980 3878
rect 51000 3398 51028 309742
rect 57256 180810 57284 405690
rect 237378 403064 237434 403073
rect 237378 402999 237380 403008
rect 237432 402999 237434 403008
rect 237380 402970 237432 402976
rect 237378 399256 237434 399265
rect 237378 399191 237434 399200
rect 237392 398886 237420 399191
rect 237380 398880 237432 398886
rect 237380 398822 237432 398828
rect 237378 396128 237434 396137
rect 237378 396063 237380 396072
rect 237432 396063 237434 396072
rect 237380 396034 237432 396040
rect 237378 390552 237434 390561
rect 237378 390487 237380 390496
rect 237432 390487 237434 390496
rect 237380 390458 237432 390464
rect 237380 387796 237432 387802
rect 237380 387738 237432 387744
rect 237392 387705 237420 387738
rect 237378 387696 237434 387705
rect 237378 387631 237434 387640
rect 237380 385008 237432 385014
rect 237378 384976 237380 384985
rect 237432 384976 237434 384985
rect 237378 384911 237434 384920
rect 237380 382220 237432 382226
rect 237380 382162 237432 382168
rect 237392 381857 237420 382162
rect 237378 381848 237434 381857
rect 237378 381783 237434 381792
rect 237380 378140 237432 378146
rect 237380 378082 237432 378088
rect 237392 378049 237420 378082
rect 237378 378040 237434 378049
rect 237378 377975 237434 377984
rect 237380 375352 237432 375358
rect 237378 375320 237380 375329
rect 237432 375320 237434 375329
rect 237378 375255 237434 375264
rect 237378 371512 237434 371521
rect 237378 371447 237434 371456
rect 237392 371278 237420 371447
rect 237380 371272 237432 371278
rect 237380 371214 237432 371220
rect 237378 365800 237434 365809
rect 237378 365735 237380 365744
rect 237432 365735 237434 365744
rect 237380 365706 237432 365712
rect 237378 358864 237434 358873
rect 237378 358799 237380 358808
rect 237432 358799 237434 358808
rect 237380 358770 237432 358776
rect 237378 352608 237434 352617
rect 237378 352543 237434 352552
rect 237392 351966 237420 352543
rect 237380 351960 237432 351966
rect 237380 351902 237432 351908
rect 237380 347744 237432 347750
rect 237378 347712 237380 347721
rect 237432 347712 237434 347721
rect 237378 347647 237434 347656
rect 237380 345024 237432 345030
rect 237380 344966 237432 344972
rect 237392 344593 237420 344966
rect 237378 344584 237434 344593
rect 237378 344519 237434 344528
rect 237380 340876 237432 340882
rect 237380 340818 237432 340824
rect 237392 340785 237420 340818
rect 237378 340776 237434 340785
rect 237378 340711 237434 340720
rect 237380 338088 237432 338094
rect 237378 338056 237380 338065
rect 237432 338056 237434 338065
rect 237378 337991 237434 338000
rect 237380 335300 237432 335306
rect 237380 335242 237432 335248
rect 237392 335209 237420 335242
rect 237378 335200 237434 335209
rect 237378 335135 237434 335144
rect 237380 332580 237432 332586
rect 237380 332522 237432 332528
rect 237392 332217 237420 332522
rect 237378 332208 237434 332217
rect 237378 332143 237434 332152
rect 229744 328092 229796 328098
rect 229744 328034 229796 328040
rect 122748 327752 122800 327758
rect 122748 327694 122800 327700
rect 104808 313948 104860 313954
rect 104808 313890 104860 313896
rect 86868 312588 86920 312594
rect 86868 312530 86920 312536
rect 57888 311160 57940 311166
rect 57888 311102 57940 311108
rect 57244 180804 57296 180810
rect 57244 180746 57296 180752
rect 55128 13116 55180 13122
rect 55128 13058 55180 13064
rect 55140 3398 55168 13058
rect 57900 6914 57928 311102
rect 62028 278044 62080 278050
rect 62028 277986 62080 277992
rect 57624 6886 57928 6914
rect 50528 3392 50580 3398
rect 50528 3334 50580 3340
rect 50988 3392 51040 3398
rect 50988 3334 51040 3340
rect 54024 3392 54076 3398
rect 54024 3334 54076 3340
rect 55128 3392 55180 3398
rect 55128 3334 55180 3340
rect 50540 480 50568 3334
rect 54036 480 54064 3334
rect 57624 480 57652 6886
rect 62040 3398 62068 277986
rect 64788 276684 64840 276690
rect 64788 276626 64840 276632
rect 61200 3392 61252 3398
rect 61200 3334 61252 3340
rect 62028 3392 62080 3398
rect 62028 3334 62080 3340
rect 61212 480 61240 3334
rect 64800 480 64828 276626
rect 73068 275324 73120 275330
rect 73068 275266 73120 275272
rect 68928 40724 68980 40730
rect 68928 40666 68980 40672
rect 68940 3398 68968 40666
rect 73080 3398 73108 275266
rect 75828 273964 75880 273970
rect 75828 273906 75880 273912
rect 75840 6914 75868 273906
rect 82728 272536 82780 272542
rect 82728 272478 82780 272484
rect 79968 44872 80020 44878
rect 79968 44814 80020 44820
rect 75472 6886 75868 6914
rect 68284 3392 68336 3398
rect 68284 3334 68336 3340
rect 68928 3392 68980 3398
rect 68928 3334 68980 3340
rect 71872 3392 71924 3398
rect 71872 3334 71924 3340
rect 73068 3392 73120 3398
rect 73068 3334 73120 3340
rect 68296 480 68324 3334
rect 71884 480 71912 3334
rect 75472 480 75500 6886
rect 79980 3398 80008 44814
rect 82740 6914 82768 272478
rect 82648 6886 82768 6914
rect 79048 3392 79100 3398
rect 79048 3334 79100 3340
rect 79968 3392 80020 3398
rect 79968 3334 80020 3340
rect 79060 480 79088 3334
rect 82648 480 82676 6886
rect 86880 2922 86908 312530
rect 93768 289128 93820 289134
rect 93768 289070 93820 289076
rect 91008 271176 91060 271182
rect 91008 271118 91060 271124
rect 91020 3398 91048 271118
rect 93780 3398 93808 289070
rect 97908 269816 97960 269822
rect 97908 269758 97960 269764
rect 97920 3398 97948 269758
rect 100668 46232 100720 46238
rect 100668 46174 100720 46180
rect 100680 6914 100708 46174
rect 100496 6886 100708 6914
rect 89720 3392 89772 3398
rect 89720 3334 89772 3340
rect 91008 3392 91060 3398
rect 91008 3334 91060 3340
rect 93308 3392 93360 3398
rect 93308 3334 93360 3340
rect 93768 3392 93820 3398
rect 93768 3334 93820 3340
rect 96896 3392 96948 3398
rect 96896 3334 96948 3340
rect 97908 3392 97960 3398
rect 97908 3334 97960 3340
rect 86132 2916 86184 2922
rect 86132 2858 86184 2864
rect 86868 2916 86920 2922
rect 86868 2858 86920 2864
rect 86144 480 86172 2858
rect 89732 480 89760 3334
rect 93320 480 93348 3334
rect 96908 480 96936 3334
rect 100496 480 100524 6886
rect 104820 3398 104848 313890
rect 107568 268388 107620 268394
rect 107568 268330 107620 268336
rect 103980 3392 104032 3398
rect 103980 3334 104032 3340
rect 104808 3392 104860 3398
rect 104808 3334 104860 3340
rect 103992 480 104020 3334
rect 107580 480 107608 268330
rect 114744 4072 114796 4078
rect 114744 4014 114796 4020
rect 111156 4004 111208 4010
rect 111156 3946 111208 3952
rect 111168 480 111196 3946
rect 114756 480 114784 4014
rect 118240 3392 118292 3398
rect 118240 3334 118292 3340
rect 118252 480 118280 3334
rect 122760 3330 122788 327694
rect 219348 326460 219400 326466
rect 219348 326402 219400 326408
rect 126888 326392 126940 326398
rect 126888 326334 126940 326340
rect 126900 6914 126928 326334
rect 162768 324964 162820 324970
rect 162768 324906 162820 324912
rect 133788 307080 133840 307086
rect 133788 307022 133840 307028
rect 132408 294636 132460 294642
rect 132408 294578 132460 294584
rect 131028 11756 131080 11762
rect 131028 11698 131080 11704
rect 126624 6886 126928 6914
rect 121828 3324 121880 3330
rect 121828 3266 121880 3272
rect 122748 3324 122800 3330
rect 122748 3266 122800 3272
rect 125416 3324 125468 3330
rect 125416 3266 125468 3272
rect 121840 480 121868 3266
rect 125428 480 125456 3266
rect 126624 480 126652 6886
rect 131040 3398 131068 11698
rect 130200 3392 130252 3398
rect 130200 3334 130252 3340
rect 131028 3392 131080 3398
rect 131028 3334 131080 3340
rect 130212 480 130240 3334
rect 132420 3330 132448 294578
rect 131396 3324 131448 3330
rect 131396 3266 131448 3272
rect 132408 3324 132460 3330
rect 132408 3266 132460 3272
rect 131408 480 131436 3266
rect 133800 480 133828 307022
rect 142068 305652 142120 305658
rect 142068 305594 142120 305600
rect 139308 287700 139360 287706
rect 139308 287642 139360 287648
rect 137928 29640 137980 29646
rect 137928 29582 137980 29588
rect 135168 26920 135220 26926
rect 135168 26862 135220 26868
rect 135180 6914 135208 26862
rect 134904 6886 135208 6914
rect 134904 480 134932 6886
rect 137940 3330 137968 29582
rect 139320 3330 139348 287642
rect 141976 286340 142028 286346
rect 141976 286282 142028 286288
rect 137284 3324 137336 3330
rect 137284 3266 137336 3272
rect 137928 3324 137980 3330
rect 137928 3266 137980 3272
rect 138480 3324 138532 3330
rect 138480 3266 138532 3272
rect 139308 3324 139360 3330
rect 139308 3266 139360 3272
rect 140872 3324 140924 3330
rect 140872 3266 140924 3272
rect 137296 480 137324 3266
rect 138492 480 138520 3266
rect 140884 480 140912 3266
rect 141988 1578 142016 286282
rect 142080 3330 142108 305594
rect 144828 304292 144880 304298
rect 144828 304234 144880 304240
rect 144840 6914 144868 304234
rect 151728 302932 151780 302938
rect 151728 302874 151780 302880
rect 146208 284980 146260 284986
rect 146208 284922 146260 284928
rect 144472 6886 144868 6914
rect 142068 3324 142120 3330
rect 142068 3266 142120 3272
rect 141988 1550 142108 1578
rect 142080 480 142108 1550
rect 144472 480 144500 6886
rect 146220 3330 146248 284922
rect 150348 283620 150400 283626
rect 150348 283562 150400 283568
rect 148968 14476 149020 14482
rect 148968 14418 149020 14424
rect 148980 3330 149008 14418
rect 150360 3330 150388 283562
rect 151740 6914 151768 302874
rect 160008 301504 160060 301510
rect 160008 301446 160060 301452
rect 159916 42084 159968 42090
rect 159916 42026 159968 42032
rect 153108 37936 153160 37942
rect 153108 37878 153160 37884
rect 153120 6914 153148 37878
rect 155868 17264 155920 17270
rect 155868 17206 155920 17212
rect 151556 6886 151768 6914
rect 152752 6886 153148 6914
rect 145656 3324 145708 3330
rect 145656 3266 145708 3272
rect 146208 3324 146260 3330
rect 146208 3266 146260 3272
rect 148048 3324 148100 3330
rect 148048 3266 148100 3272
rect 148968 3324 149020 3330
rect 148968 3266 149020 3272
rect 149244 3324 149296 3330
rect 149244 3266 149296 3272
rect 150348 3324 150400 3330
rect 150348 3266 150400 3272
rect 145668 480 145696 3266
rect 148060 480 148088 3266
rect 149256 480 149284 3266
rect 151556 480 151584 6886
rect 152752 480 152780 6886
rect 155880 3330 155908 17206
rect 157248 10328 157300 10334
rect 157248 10270 157300 10276
rect 157260 3330 157288 10270
rect 155132 3324 155184 3330
rect 155132 3266 155184 3272
rect 155868 3324 155920 3330
rect 155868 3266 155920 3272
rect 156328 3324 156380 3330
rect 156328 3266 156380 3272
rect 157248 3324 157300 3330
rect 157248 3266 157300 3272
rect 158720 3324 158772 3330
rect 158720 3266 158772 3272
rect 155144 480 155172 3266
rect 156340 480 156368 3266
rect 158732 480 158760 3266
rect 159928 480 159956 42026
rect 160020 3330 160048 301446
rect 162780 3330 162808 324906
rect 169668 322244 169720 322250
rect 169668 322186 169720 322192
rect 168288 300144 168340 300150
rect 168288 300086 168340 300092
rect 164148 19984 164200 19990
rect 164148 19926 164200 19932
rect 164160 3330 164188 19926
rect 165896 4820 165948 4826
rect 165896 4762 165948 4768
rect 160008 3324 160060 3330
rect 160008 3266 160060 3272
rect 162308 3324 162360 3330
rect 162308 3266 162360 3272
rect 162768 3324 162820 3330
rect 162768 3266 162820 3272
rect 163504 3324 163556 3330
rect 163504 3266 163556 3272
rect 164148 3324 164200 3330
rect 164148 3266 164200 3272
rect 162320 480 162348 3266
rect 163516 480 163544 3266
rect 165908 480 165936 4762
rect 168300 3330 168328 300086
rect 169680 6914 169708 322186
rect 176568 320884 176620 320890
rect 176568 320826 176620 320832
rect 175188 21412 175240 21418
rect 175188 21354 175240 21360
rect 171048 18624 171100 18630
rect 171048 18566 171100 18572
rect 169404 6886 169708 6914
rect 167092 3324 167144 3330
rect 167092 3266 167144 3272
rect 168288 3324 168340 3330
rect 168288 3266 168340 3272
rect 167104 480 167132 3266
rect 169404 480 169432 6886
rect 171060 3330 171088 18566
rect 172980 6180 173032 6186
rect 172980 6122 173032 6128
rect 170588 3324 170640 3330
rect 170588 3266 170640 3272
rect 171048 3324 171100 3330
rect 171048 3266 171100 3272
rect 170600 480 170628 3266
rect 172992 480 173020 6122
rect 175200 3330 175228 21354
rect 174176 3324 174228 3330
rect 174176 3266 174228 3272
rect 175188 3324 175240 3330
rect 175188 3266 175240 3272
rect 174188 480 174216 3266
rect 176580 480 176608 320826
rect 180708 319456 180760 319462
rect 180708 319398 180760 319404
rect 177948 298784 178000 298790
rect 177948 298726 178000 298732
rect 177960 6914 177988 298726
rect 177776 6886 177988 6914
rect 177776 480 177804 6886
rect 180720 3330 180748 319398
rect 187608 318096 187660 318102
rect 187608 318038 187660 318044
rect 184848 25560 184900 25566
rect 184848 25502 184900 25508
rect 182088 22772 182140 22778
rect 182088 22714 182140 22720
rect 182100 3330 182128 22714
rect 183744 8968 183796 8974
rect 183744 8910 183796 8916
rect 180156 3324 180208 3330
rect 180156 3266 180208 3272
rect 180708 3324 180760 3330
rect 180708 3266 180760 3272
rect 181352 3324 181404 3330
rect 181352 3266 181404 3272
rect 182088 3324 182140 3330
rect 182088 3266 182140 3272
rect 180168 480 180196 3266
rect 181364 480 181392 3266
rect 183756 480 183784 8910
rect 184860 480 184888 25502
rect 187620 6914 187648 318038
rect 194508 316736 194560 316742
rect 194508 316678 194560 316684
rect 193128 297424 193180 297430
rect 193128 297366 193180 297372
rect 188988 24132 189040 24138
rect 188988 24074 189040 24080
rect 187252 6886 187648 6914
rect 187252 480 187280 6886
rect 189000 3194 189028 24074
rect 191748 15904 191800 15910
rect 191748 15846 191800 15852
rect 191760 3330 191788 15846
rect 193140 3330 193168 297366
rect 194520 6914 194548 316678
rect 198648 315308 198700 315314
rect 198648 315250 198700 315256
rect 195888 295996 195940 296002
rect 195888 295938 195940 295944
rect 195900 6914 195928 295938
rect 194428 6886 194548 6914
rect 195624 6886 195928 6914
rect 190828 3324 190880 3330
rect 190828 3266 190880 3272
rect 191748 3324 191800 3330
rect 191748 3266 191800 3272
rect 192024 3324 192076 3330
rect 192024 3266 192076 3272
rect 193128 3324 193180 3330
rect 193128 3266 193180 3272
rect 188436 3188 188488 3194
rect 188436 3130 188488 3136
rect 188988 3188 189040 3194
rect 188988 3130 189040 3136
rect 188448 480 188476 3130
rect 190840 480 190868 3266
rect 192036 480 192064 3266
rect 194428 480 194456 6886
rect 195624 480 195652 6886
rect 198660 3330 198688 315250
rect 205548 314016 205600 314022
rect 205548 313958 205600 313964
rect 202788 293276 202840 293282
rect 202788 293218 202840 293224
rect 202696 91792 202748 91798
rect 202696 91734 202748 91740
rect 200028 28280 200080 28286
rect 200028 28222 200080 28228
rect 200040 3330 200068 28222
rect 202708 6914 202736 91734
rect 202616 6886 202736 6914
rect 202616 3330 202644 6886
rect 202800 3482 202828 293218
rect 202708 3454 202828 3482
rect 198004 3324 198056 3330
rect 198004 3266 198056 3272
rect 198648 3324 198700 3330
rect 198648 3266 198700 3272
rect 199200 3324 199252 3330
rect 199200 3266 199252 3272
rect 200028 3324 200080 3330
rect 200028 3266 200080 3272
rect 201500 3324 201552 3330
rect 201500 3266 201552 3272
rect 202604 3324 202656 3330
rect 202604 3266 202656 3272
rect 198016 480 198044 3266
rect 199212 480 199240 3266
rect 201512 480 201540 3266
rect 202708 480 202736 3454
rect 205560 3330 205588 313958
rect 209688 312656 209740 312662
rect 209688 312598 209740 312604
rect 206928 32428 206980 32434
rect 206928 32370 206980 32376
rect 206940 3330 206968 32370
rect 209700 3330 209728 312598
rect 212448 311228 212500 311234
rect 212448 311170 212500 311176
rect 211068 291848 211120 291854
rect 211068 291790 211120 291796
rect 211080 3330 211108 291790
rect 212460 6914 212488 311170
rect 216588 309868 216640 309874
rect 216588 309810 216640 309816
rect 213828 290488 213880 290494
rect 213828 290430 213880 290436
rect 213840 6914 213868 290430
rect 212276 6886 212488 6914
rect 213472 6886 213868 6914
rect 205088 3324 205140 3330
rect 205088 3266 205140 3272
rect 205548 3324 205600 3330
rect 205548 3266 205600 3272
rect 206284 3324 206336 3330
rect 206284 3266 206336 3272
rect 206928 3324 206980 3330
rect 206928 3266 206980 3272
rect 208676 3324 208728 3330
rect 208676 3266 208728 3272
rect 209688 3324 209740 3330
rect 209688 3266 209740 3272
rect 209872 3324 209924 3330
rect 209872 3266 209924 3272
rect 211068 3324 211120 3330
rect 211068 3266 211120 3272
rect 205100 480 205128 3266
rect 206296 480 206324 3266
rect 208688 480 208716 3266
rect 209884 480 209912 3266
rect 212276 480 212304 6886
rect 213472 480 213500 6886
rect 216600 3330 216628 309810
rect 217968 31068 218020 31074
rect 217968 31010 218020 31016
rect 217980 3330 218008 31010
rect 215852 3324 215904 3330
rect 215852 3266 215904 3272
rect 216588 3324 216640 3330
rect 216588 3266 216640 3272
rect 217048 3324 217100 3330
rect 217048 3266 217100 3272
rect 217968 3324 218020 3330
rect 217968 3266 218020 3272
rect 215864 480 215892 3266
rect 217060 480 217088 3266
rect 219360 480 219388 326402
rect 227628 323604 227680 323610
rect 227628 323546 227680 323552
rect 223488 308508 223540 308514
rect 223488 308450 223540 308456
rect 220728 33788 220780 33794
rect 220728 33730 220780 33736
rect 220740 6914 220768 33730
rect 220556 6886 220768 6914
rect 220556 480 220584 6886
rect 223500 3330 223528 308450
rect 224868 35216 224920 35222
rect 224868 35158 224920 35164
rect 224880 3330 224908 35158
rect 227640 3330 227668 323546
rect 229008 289196 229060 289202
rect 229008 289138 229060 289144
rect 229020 3330 229048 289138
rect 229756 13122 229784 328034
rect 236644 328024 236696 328030
rect 236644 327966 236696 327972
rect 231124 327956 231176 327962
rect 231124 327898 231176 327904
rect 229744 13116 229796 13122
rect 229744 13058 229796 13064
rect 230112 13116 230164 13122
rect 230112 13058 230164 13064
rect 222936 3324 222988 3330
rect 222936 3266 222988 3272
rect 223488 3324 223540 3330
rect 223488 3266 223540 3272
rect 224132 3324 224184 3330
rect 224132 3266 224184 3272
rect 224868 3324 224920 3330
rect 224868 3266 224920 3272
rect 226524 3324 226576 3330
rect 226524 3266 226576 3272
rect 227628 3324 227680 3330
rect 227628 3266 227680 3272
rect 227720 3324 227772 3330
rect 227720 3266 227772 3272
rect 229008 3324 229060 3330
rect 229008 3266 229060 3272
rect 222948 480 222976 3266
rect 224144 480 224172 3266
rect 226536 480 226564 3266
rect 227732 480 227760 3266
rect 230124 480 230152 13058
rect 231136 11762 231164 327898
rect 233884 327888 233936 327894
rect 233884 327830 233936 327836
rect 232504 327820 232556 327826
rect 232504 327762 232556 327768
rect 231768 322312 231820 322318
rect 231768 322254 231820 322260
rect 231124 11756 231176 11762
rect 231124 11698 231176 11704
rect 231780 3330 231808 322254
rect 232516 8974 232544 327762
rect 232504 8968 232556 8974
rect 232504 8910 232556 8916
rect 233896 6186 233924 327830
rect 235908 39364 235960 39370
rect 235908 39306 235960 39312
rect 233884 6180 233936 6186
rect 233884 6122 233936 6128
rect 233700 6112 233752 6118
rect 233700 6054 233752 6060
rect 231308 3324 231360 3330
rect 231308 3266 231360 3272
rect 231768 3324 231820 3330
rect 231768 3266 231820 3272
rect 231320 480 231348 3266
rect 233712 480 233740 6054
rect 235920 3330 235948 39306
rect 236656 4826 236684 327966
rect 237288 89004 237340 89010
rect 237288 88946 237340 88952
rect 237300 6914 237328 88946
rect 238036 8294 238064 418231
rect 321836 416764 321888 416770
rect 321836 416706 321888 416712
rect 321848 416401 321876 416706
rect 321834 416392 321890 416401
rect 321834 416327 321890 416336
rect 322204 413976 322256 413982
rect 322204 413918 322256 413924
rect 322216 413545 322244 413918
rect 322202 413536 322258 413545
rect 322202 413471 322258 413480
rect 238114 411632 238170 411641
rect 238114 411567 238170 411576
rect 238128 93838 238156 411567
rect 380176 411262 380204 509254
rect 384316 413982 384344 556174
rect 391204 545148 391256 545154
rect 391204 545090 391256 545096
rect 388444 498228 388496 498234
rect 388444 498170 388496 498176
rect 384304 413976 384356 413982
rect 384304 413918 384356 413924
rect 322204 411256 322256 411262
rect 322204 411198 322256 411204
rect 380164 411256 380216 411262
rect 380164 411198 380216 411204
rect 322216 410825 322244 411198
rect 322202 410816 322258 410825
rect 322202 410751 322258 410760
rect 322020 408468 322072 408474
rect 322020 408410 322072 408416
rect 322032 408105 322060 408410
rect 322018 408096 322074 408105
rect 322018 408031 322074 408040
rect 321836 405680 321888 405686
rect 321836 405622 321888 405628
rect 321848 405385 321876 405622
rect 321834 405376 321890 405385
rect 321834 405311 321890 405320
rect 322110 401704 322166 401713
rect 322110 401639 322166 401648
rect 238298 393408 238354 393417
rect 238298 393343 238354 393352
rect 238206 368520 238262 368529
rect 238206 368455 238262 368464
rect 238116 93832 238168 93838
rect 238116 93774 238168 93780
rect 238220 64870 238248 368455
rect 238312 367062 238340 393343
rect 322124 393314 322152 401639
rect 322754 398984 322810 398993
rect 322754 398919 322810 398928
rect 322202 396536 322258 396545
rect 322202 396471 322258 396480
rect 322216 396098 322244 396471
rect 322204 396092 322256 396098
rect 322204 396034 322256 396040
rect 322480 394664 322532 394670
rect 322480 394606 322532 394612
rect 322492 394369 322520 394606
rect 322478 394360 322534 394369
rect 322478 394295 322534 394304
rect 322124 393286 322244 393314
rect 321834 371784 321890 371793
rect 321834 371719 321890 371728
rect 321848 371278 321876 371719
rect 321836 371272 321888 371278
rect 321836 371214 321888 371220
rect 322216 369850 322244 393286
rect 322480 391944 322532 391950
rect 322480 391886 322532 391892
rect 322492 391649 322520 391886
rect 322478 391640 322534 391649
rect 322478 391575 322534 391584
rect 322480 389156 322532 389162
rect 322480 389098 322532 389104
rect 322492 388929 322520 389098
rect 322478 388920 322534 388929
rect 322478 388855 322534 388864
rect 322480 386368 322532 386374
rect 322480 386310 322532 386316
rect 322492 386209 322520 386310
rect 322478 386200 322534 386209
rect 322478 386135 322534 386144
rect 322480 383648 322532 383654
rect 322480 383590 322532 383596
rect 322492 383489 322520 383590
rect 322478 383480 322534 383489
rect 322478 383415 322534 383424
rect 322480 380860 322532 380866
rect 322480 380802 322532 380808
rect 322492 380769 322520 380802
rect 322478 380760 322534 380769
rect 322478 380695 322534 380704
rect 322480 378140 322532 378146
rect 322480 378082 322532 378088
rect 322492 378049 322520 378082
rect 322478 378040 322534 378049
rect 322478 377975 322534 377984
rect 322294 374504 322350 374513
rect 322294 374439 322350 374448
rect 322204 369844 322256 369850
rect 322204 369786 322256 369792
rect 238300 367056 238352 367062
rect 238300 366998 238352 367004
rect 321834 363488 321890 363497
rect 321834 363423 321890 363432
rect 321848 362982 321876 363423
rect 321836 362976 321888 362982
rect 321836 362918 321888 362924
rect 238298 361992 238354 362001
rect 238298 361927 238354 361936
rect 238312 151774 238340 361927
rect 321834 360768 321890 360777
rect 321834 360703 321890 360712
rect 321848 360262 321876 360703
rect 321836 360256 321888 360262
rect 321836 360198 321888 360204
rect 322308 358766 322336 374439
rect 322662 368928 322718 368937
rect 322662 368863 322718 368872
rect 322570 366208 322626 366217
rect 322570 366143 322626 366152
rect 322296 358760 322348 358766
rect 322296 358702 322348 358708
rect 322478 358048 322534 358057
rect 322478 357983 322534 357992
rect 238390 356144 238446 356153
rect 238390 356079 238446 356088
rect 238404 237386 238432 356079
rect 321650 355600 321706 355609
rect 321650 355535 321706 355544
rect 321664 355162 321692 355535
rect 321652 355156 321704 355162
rect 321652 355098 321704 355104
rect 322386 352608 322442 352617
rect 322386 352543 322442 352552
rect 322018 349888 322074 349897
rect 322018 349823 322074 349832
rect 238482 349480 238538 349489
rect 238482 349415 238538 349424
rect 238496 324290 238524 349415
rect 322032 349178 322060 349823
rect 322020 349172 322072 349178
rect 322020 349114 322072 349120
rect 322018 347168 322074 347177
rect 322018 347103 322074 347112
rect 322032 346458 322060 347103
rect 322020 346452 322072 346458
rect 322020 346394 322072 346400
rect 322294 345128 322350 345137
rect 322294 345063 322296 345072
rect 322348 345063 322350 345072
rect 322296 345034 322348 345040
rect 322202 342272 322258 342281
rect 322202 342207 322258 342216
rect 322216 339402 322244 342207
rect 322294 339552 322350 339561
rect 322294 339487 322296 339496
rect 322348 339487 322350 339496
rect 322296 339458 322348 339464
rect 322216 339374 322336 339402
rect 322202 336832 322258 336841
rect 322202 336767 322258 336776
rect 322110 334112 322166 334121
rect 322110 334047 322166 334056
rect 322124 334014 322152 334047
rect 322112 334008 322164 334014
rect 322112 333950 322164 333956
rect 322110 331392 322166 331401
rect 322110 331327 322166 331336
rect 322124 331294 322152 331327
rect 322112 331288 322164 331294
rect 322112 331230 322164 331236
rect 240258 330126 240364 330154
rect 243018 330126 243124 330154
rect 247158 330126 247356 330154
rect 251206 330126 251312 330154
rect 258106 330126 258212 330154
rect 271078 330126 271368 330154
rect 271538 330126 271736 330154
rect 271906 330126 272104 330154
rect 272274 330126 272564 330154
rect 272734 330126 272932 330154
rect 273562 330126 273760 330154
rect 273930 330126 274128 330154
rect 274298 330126 274404 330154
rect 274758 330126 274956 330154
rect 275586 330126 275784 330154
rect 276414 330126 276612 330154
rect 276782 330126 276980 330154
rect 277150 330126 277256 330154
rect 278806 330126 279004 330154
rect 279174 330126 279464 330154
rect 279634 330126 279832 330154
rect 280462 330126 280660 330154
rect 280830 330126 281120 330154
rect 281290 330126 281488 330154
rect 285706 330126 285812 330154
rect 292606 330126 292712 330154
rect 299506 330126 299612 330154
rect 301162 330126 301360 330154
rect 301530 330126 301820 330154
rect 302358 330126 302648 330154
rect 302818 330126 303016 330154
rect 303186 330126 303384 330154
rect 304014 330126 304212 330154
rect 304382 330126 304672 330154
rect 305210 330126 305500 330154
rect 305670 330126 305868 330154
rect 306038 330126 306236 330154
rect 306406 330126 306696 330154
rect 306866 330126 307064 330154
rect 307234 330126 307524 330154
rect 308062 330126 308260 330154
rect 308430 330126 308720 330154
rect 308890 330126 308996 330154
rect 309258 330126 309364 330154
rect 310086 330126 310284 330154
rect 310546 330126 310652 330154
rect 310914 330126 311112 330154
rect 311282 330126 311480 330154
rect 312110 330126 312400 330154
rect 312570 330126 312768 330154
rect 312938 330126 313136 330154
rect 313306 330126 313412 330154
rect 314134 330126 314424 330154
rect 314962 330126 315252 330154
rect 315422 330126 315620 330154
rect 315790 330126 315896 330154
rect 316158 330126 316448 330154
rect 316618 330126 316816 330154
rect 316986 330126 317276 330154
rect 317446 330126 317644 330154
rect 317814 330126 318012 330154
rect 318182 330126 318472 330154
rect 318642 330126 318748 330154
rect 319010 330126 319300 330154
rect 319470 330126 319668 330154
rect 319838 330126 320128 330154
rect 239404 328160 239456 328166
rect 239404 328102 239456 328108
rect 239416 326398 239444 328102
rect 239404 326392 239456 326398
rect 239404 326334 239456 326340
rect 238484 324284 238536 324290
rect 238484 324226 238536 324232
rect 240336 282198 240364 330126
rect 240520 329990 240626 330018
rect 240704 329990 240994 330018
rect 241072 329990 241454 330018
rect 241624 329990 241822 330018
rect 241900 329990 242282 330018
rect 242360 329990 242650 330018
rect 240416 325780 240468 325786
rect 240416 325722 240468 325728
rect 240324 282192 240376 282198
rect 240324 282134 240376 282140
rect 238392 237380 238444 237386
rect 238392 237322 238444 237328
rect 238300 151768 238352 151774
rect 238300 151710 238352 151716
rect 238208 64864 238260 64870
rect 238208 64806 238260 64812
rect 238668 36576 238720 36582
rect 238668 36518 238720 36524
rect 238024 8288 238076 8294
rect 238024 8230 238076 8236
rect 238680 6914 238708 36518
rect 237208 6886 237328 6914
rect 238404 6886 238708 6914
rect 236644 4820 236696 4826
rect 236644 4762 236696 4768
rect 234804 3324 234856 3330
rect 234804 3266 234856 3272
rect 235908 3324 235960 3330
rect 235908 3266 235960 3272
rect 234816 480 234844 3266
rect 237208 480 237236 6886
rect 238404 480 238432 6886
rect 240428 3398 240456 325722
rect 240520 280838 240548 329990
rect 240704 327758 240732 329990
rect 240692 327752 240744 327758
rect 240692 327694 240744 327700
rect 241072 325786 241100 329990
rect 241060 325780 241112 325786
rect 241060 325722 241112 325728
rect 241520 325780 241572 325786
rect 241520 325722 241572 325728
rect 240508 280832 240560 280838
rect 240508 280774 240560 280780
rect 241532 271182 241560 325722
rect 241624 308446 241652 329990
rect 241900 312594 241928 329990
rect 242360 325786 242388 329990
rect 242348 325780 242400 325786
rect 242348 325722 242400 325728
rect 241888 312588 241940 312594
rect 241888 312530 241940 312536
rect 241612 308440 241664 308446
rect 241612 308382 241664 308388
rect 243096 289134 243124 330126
rect 243372 329990 243478 330018
rect 243556 329990 243846 330018
rect 244246 329990 244306 330018
rect 244476 329990 244674 330018
rect 244752 329990 245042 330018
rect 245120 329990 245502 330018
rect 245764 329990 245870 330018
rect 245948 329990 246330 330018
rect 246408 329990 246698 330018
rect 243372 325650 243400 329990
rect 243360 325644 243412 325650
rect 243360 325586 243412 325592
rect 243268 325440 243320 325446
rect 243268 325382 243320 325388
rect 243176 323672 243228 323678
rect 243176 323614 243228 323620
rect 243084 289128 243136 289134
rect 243084 289070 243136 289076
rect 241520 271176 241572 271182
rect 241520 271118 241572 271124
rect 243188 46238 243216 323614
rect 243280 269822 243308 325382
rect 243556 323678 243584 329990
rect 244246 329882 244274 329990
rect 244246 329854 244320 329882
rect 243544 323672 243596 323678
rect 243544 323614 243596 323620
rect 244292 313954 244320 329854
rect 244372 325780 244424 325786
rect 244372 325722 244424 325728
rect 244280 313948 244332 313954
rect 244280 313890 244332 313896
rect 243268 269816 243320 269822
rect 243268 269758 243320 269764
rect 243176 46232 243228 46238
rect 243176 46174 243228 46180
rect 242808 11756 242860 11762
rect 242808 11698 242860 11704
rect 240784 4888 240836 4894
rect 240784 4830 240836 4836
rect 240416 3392 240468 3398
rect 240416 3334 240468 3340
rect 240796 480 240824 4830
rect 242820 3398 242848 11698
rect 244384 4010 244412 325722
rect 244476 268394 244504 329990
rect 244752 325786 244780 329990
rect 244740 325780 244792 325786
rect 244740 325722 244792 325728
rect 245120 316034 245148 329990
rect 245764 321554 245792 329990
rect 245764 321526 245884 321554
rect 244752 316006 245148 316034
rect 244464 268388 244516 268394
rect 244464 268330 244516 268336
rect 244464 7676 244516 7682
rect 244464 7618 244516 7624
rect 244372 4004 244424 4010
rect 244372 3946 244424 3952
rect 244476 3482 244504 7618
rect 244752 4078 244780 316006
rect 245568 4820 245620 4826
rect 245568 4762 245620 4768
rect 244740 4072 244792 4078
rect 244740 4014 244792 4020
rect 244384 3454 244504 3482
rect 241980 3392 242032 3398
rect 241980 3334 242032 3340
rect 242808 3392 242860 3398
rect 242808 3334 242860 3340
rect 241992 480 242020 3334
rect 244384 480 244412 3454
rect 245580 480 245608 4762
rect 245856 4146 245884 321526
rect 245948 309806 245976 329990
rect 246408 328098 246436 329990
rect 246396 328092 246448 328098
rect 246396 328034 246448 328040
rect 247328 325922 247356 330126
rect 247420 329990 247526 330018
rect 247696 329990 247894 330018
rect 248064 329990 248354 330018
rect 248616 329990 248722 330018
rect 248800 329990 249182 330018
rect 249260 329990 249550 330018
rect 249812 329990 249918 330018
rect 249996 329990 250378 330018
rect 250456 329990 250746 330018
rect 247316 325916 247368 325922
rect 247316 325858 247368 325864
rect 247316 325712 247368 325718
rect 247316 325654 247368 325660
rect 247224 323672 247276 323678
rect 247224 323614 247276 323620
rect 245936 309800 245988 309806
rect 245936 309742 245988 309748
rect 247236 278050 247264 323614
rect 247328 311166 247356 325654
rect 247420 323678 247448 329990
rect 247592 325780 247644 325786
rect 247592 325722 247644 325728
rect 247408 323672 247460 323678
rect 247408 323614 247460 323620
rect 247316 311160 247368 311166
rect 247316 311102 247368 311108
rect 247224 278044 247276 278050
rect 247224 277986 247276 277992
rect 247604 40730 247632 325722
rect 247696 276690 247724 329990
rect 248064 325786 248092 329990
rect 248616 325922 248644 329990
rect 248800 328454 248828 329990
rect 248708 328426 248828 328454
rect 248604 325916 248656 325922
rect 248604 325858 248656 325864
rect 248052 325780 248104 325786
rect 248052 325722 248104 325728
rect 248420 325780 248472 325786
rect 248420 325722 248472 325728
rect 247684 276684 247736 276690
rect 247684 276626 247736 276632
rect 248432 44878 248460 325722
rect 248708 323762 248736 328426
rect 249260 325786 249288 329990
rect 249248 325780 249300 325786
rect 249248 325722 249300 325728
rect 248524 323734 248736 323762
rect 248524 273970 248552 323734
rect 248604 323672 248656 323678
rect 248604 323614 248656 323620
rect 248616 275330 248644 323614
rect 249812 321554 249840 329990
rect 249812 321526 249932 321554
rect 248604 275324 248656 275330
rect 248604 275266 248656 275272
rect 248512 273964 248564 273970
rect 248512 273906 248564 273912
rect 249904 272542 249932 321526
rect 249996 279478 250024 329990
rect 250456 316034 250484 329990
rect 250088 316006 250484 316034
rect 249984 279472 250036 279478
rect 249984 279414 250036 279420
rect 249892 272536 249944 272542
rect 249892 272478 249944 272484
rect 248420 44872 248472 44878
rect 248420 44814 248472 44820
rect 250088 43450 250116 316006
rect 250076 43444 250128 43450
rect 250076 43386 250128 43392
rect 247592 40724 247644 40730
rect 247592 40666 247644 40672
rect 249708 29708 249760 29714
rect 249708 29650 249760 29656
rect 247960 9036 248012 9042
rect 247960 8978 248012 8984
rect 245844 4140 245896 4146
rect 245844 4082 245896 4088
rect 247972 480 248000 8978
rect 249720 3534 249748 29650
rect 249156 3528 249208 3534
rect 249156 3470 249208 3476
rect 249708 3528 249760 3534
rect 249708 3470 249760 3476
rect 249168 480 249196 3470
rect 251284 3466 251312 330126
rect 251376 329990 251574 330018
rect 251744 329990 252034 330018
rect 252112 329990 252402 330018
rect 252664 329990 252770 330018
rect 252848 329990 253230 330018
rect 253308 329990 253598 330018
rect 253952 329990 254058 330018
rect 254136 329990 254426 330018
rect 254504 329990 254794 330018
rect 254872 329990 255254 330018
rect 255332 329990 255622 330018
rect 255700 329990 256082 330018
rect 256160 329990 256450 330018
rect 256712 329990 256910 330018
rect 257172 329990 257278 330018
rect 257356 329990 257646 330018
rect 251376 3602 251404 329990
rect 251640 325780 251692 325786
rect 251640 325722 251692 325728
rect 251456 6248 251508 6254
rect 251456 6190 251508 6196
rect 251364 3596 251416 3602
rect 251364 3538 251416 3544
rect 251272 3460 251324 3466
rect 251272 3402 251324 3408
rect 251468 480 251496 6190
rect 251652 3670 251680 325722
rect 251744 3738 251772 329990
rect 252112 325786 252140 329990
rect 252100 325780 252152 325786
rect 252100 325722 252152 325728
rect 252560 325780 252612 325786
rect 252560 325722 252612 325728
rect 252572 3874 252600 325722
rect 252664 16574 252692 329990
rect 252664 16546 252784 16574
rect 252652 7608 252704 7614
rect 252652 7550 252704 7556
rect 252560 3868 252612 3874
rect 252560 3810 252612 3816
rect 251732 3732 251784 3738
rect 251732 3674 251784 3680
rect 251640 3664 251692 3670
rect 251640 3606 251692 3612
rect 252664 480 252692 7550
rect 252756 4010 252784 16546
rect 252744 4004 252796 4010
rect 252744 3946 252796 3952
rect 252848 3806 252876 329990
rect 253308 325786 253336 329990
rect 253296 325780 253348 325786
rect 253296 325722 253348 325728
rect 253952 3942 253980 329990
rect 254136 328166 254164 329990
rect 254124 328160 254176 328166
rect 254124 328102 254176 328108
rect 254504 328098 254532 329990
rect 254492 328092 254544 328098
rect 254492 328034 254544 328040
rect 254872 325802 254900 329990
rect 255332 327162 255360 329990
rect 254504 325774 254900 325802
rect 255148 327134 255360 327162
rect 254504 307086 254532 325774
rect 255148 321554 255176 327134
rect 255700 325938 255728 329990
rect 254596 321526 255176 321554
rect 255424 325910 255728 325938
rect 254492 307080 254544 307086
rect 254492 307022 254544 307028
rect 254596 29646 254624 321526
rect 255424 305658 255452 325910
rect 256160 325802 256188 329990
rect 256712 327146 256740 329990
rect 256240 327140 256292 327146
rect 256240 327082 256292 327088
rect 256700 327140 256752 327146
rect 256700 327082 256752 327088
rect 255700 325774 256188 325802
rect 255412 305652 255464 305658
rect 255412 305594 255464 305600
rect 255700 304298 255728 325774
rect 256252 321554 256280 327082
rect 257172 325650 257200 329990
rect 257160 325644 257212 325650
rect 257160 325586 257212 325592
rect 257068 325440 257120 325446
rect 257068 325382 257120 325388
rect 255976 321526 256280 321554
rect 255688 304292 255740 304298
rect 255688 304234 255740 304240
rect 254584 29640 254636 29646
rect 254584 29582 254636 29588
rect 255228 26988 255280 26994
rect 255228 26930 255280 26936
rect 255240 6914 255268 26930
rect 255976 14482 256004 321526
rect 256976 318844 257028 318850
rect 256976 318786 257028 318792
rect 256608 304292 256660 304298
rect 256608 304234 256660 304240
rect 255964 14476 256016 14482
rect 255964 14418 256016 14424
rect 256620 6914 256648 304234
rect 256988 17270 257016 318786
rect 257080 302938 257108 325382
rect 257356 318850 257384 329990
rect 258184 321554 258212 330126
rect 258276 329990 258474 330018
rect 258552 329990 258934 330018
rect 259012 329990 259302 330018
rect 259472 329990 259670 330018
rect 259840 329990 260130 330018
rect 260208 329990 260498 330018
rect 260852 329990 260958 330018
rect 261036 329990 261326 330018
rect 261404 329990 261786 330018
rect 261864 329990 262154 330018
rect 262416 329990 262522 330018
rect 262600 329990 262982 330018
rect 263060 329990 263350 330018
rect 263612 329990 263810 330018
rect 263888 329990 264178 330018
rect 264256 329990 264546 330018
rect 264900 329990 265006 330018
rect 265084 329990 265374 330018
rect 265452 329990 265834 330018
rect 265912 329990 266202 330018
rect 266372 329990 266662 330018
rect 266740 329990 267030 330018
rect 267108 329990 267398 330018
rect 267752 329990 267858 330018
rect 267936 329990 268226 330018
rect 268304 329990 268686 330018
rect 268764 329990 269054 330018
rect 269132 329990 269422 330018
rect 269500 329990 269882 330018
rect 269960 329990 270250 330018
rect 270512 329990 270710 330018
rect 258276 324970 258304 329990
rect 258552 328030 258580 329990
rect 258540 328024 258592 328030
rect 258540 327966 258592 327972
rect 258724 327956 258776 327962
rect 258724 327898 258776 327904
rect 258356 327140 258408 327146
rect 258356 327082 258408 327088
rect 258264 324964 258316 324970
rect 258264 324906 258316 324912
rect 258092 321526 258212 321554
rect 257344 318844 257396 318850
rect 257344 318786 257396 318792
rect 257068 302932 257120 302938
rect 257068 302874 257120 302880
rect 258092 301510 258120 321526
rect 258368 320890 258396 327082
rect 258356 320884 258408 320890
rect 258356 320826 258408 320832
rect 258080 301504 258132 301510
rect 258080 301446 258132 301452
rect 256976 17264 257028 17270
rect 256976 17206 257028 17212
rect 258632 9648 258684 9654
rect 258632 9590 258684 9596
rect 255056 6886 255268 6914
rect 256252 6886 256648 6914
rect 253940 3936 253992 3942
rect 253940 3878 253992 3884
rect 252836 3800 252888 3806
rect 252836 3742 252888 3748
rect 255056 480 255084 6886
rect 256252 480 256280 6886
rect 258644 480 258672 9590
rect 258736 9042 258764 327898
rect 258816 327616 258868 327622
rect 258816 327558 258868 327564
rect 258828 26926 258856 327558
rect 259012 322250 259040 329990
rect 259472 327894 259500 329990
rect 259460 327888 259512 327894
rect 259460 327830 259512 327836
rect 259840 327146 259868 329990
rect 259828 327140 259880 327146
rect 259828 327082 259880 327088
rect 259000 322244 259052 322250
rect 259000 322186 259052 322192
rect 260208 319462 260236 329990
rect 260852 327826 260880 329990
rect 260840 327820 260892 327826
rect 260840 327762 260892 327768
rect 260196 319456 260248 319462
rect 260196 319398 260248 319404
rect 261036 318102 261064 329990
rect 261404 325938 261432 329990
rect 261128 325910 261432 325938
rect 261024 318096 261076 318102
rect 261024 318038 261076 318044
rect 260748 312588 260800 312594
rect 260748 312530 260800 312536
rect 258816 26920 258868 26926
rect 258816 26862 258868 26868
rect 258724 9036 258776 9042
rect 258724 8978 258776 8984
rect 260760 3534 260788 312530
rect 261128 15910 261156 325910
rect 261864 325802 261892 329990
rect 262036 327548 262088 327554
rect 262036 327490 262088 327496
rect 261944 327344 261996 327350
rect 261944 327286 261996 327292
rect 261404 325774 261892 325802
rect 261404 316742 261432 325774
rect 261956 324442 261984 327286
rect 261496 324414 261984 324442
rect 261392 316736 261444 316742
rect 261392 316678 261444 316684
rect 261116 15904 261168 15910
rect 261116 15846 261168 15852
rect 261496 9654 261524 324414
rect 262048 321554 262076 327490
rect 262416 326330 262444 329990
rect 262404 326324 262456 326330
rect 262404 326266 262456 326272
rect 262496 326120 262548 326126
rect 262496 326062 262548 326068
rect 262312 325712 262364 325718
rect 262312 325654 262364 325660
rect 261588 321526 262076 321554
rect 261588 312662 261616 321526
rect 262220 319048 262272 319054
rect 262220 318990 262272 318996
rect 261576 312656 261628 312662
rect 261576 312598 261628 312604
rect 262232 91798 262260 318990
rect 262324 314022 262352 325654
rect 262508 316034 262536 326062
rect 262600 319054 262628 329990
rect 262864 327684 262916 327690
rect 262864 327626 262916 327632
rect 262588 319048 262640 319054
rect 262588 318990 262640 318996
rect 262416 316006 262536 316034
rect 262416 315314 262444 316006
rect 262404 315308 262456 315314
rect 262404 315250 262456 315256
rect 262312 314016 262364 314022
rect 262312 313958 262364 313964
rect 262220 91792 262272 91798
rect 262220 91734 262272 91740
rect 261484 9648 261536 9654
rect 261484 9590 261536 9596
rect 262220 8356 262272 8362
rect 262220 8298 262272 8304
rect 259828 3528 259880 3534
rect 259828 3470 259880 3476
rect 260748 3528 260800 3534
rect 260748 3470 260800 3476
rect 259840 480 259868 3470
rect 262232 480 262260 8298
rect 262876 6186 262904 327626
rect 262956 327412 263008 327418
rect 262956 327354 263008 327360
rect 262968 311234 262996 327354
rect 263060 325718 263088 329990
rect 263612 327554 263640 329990
rect 263600 327548 263652 327554
rect 263600 327490 263652 327496
rect 263888 327418 263916 329990
rect 263876 327412 263928 327418
rect 263876 327354 263928 327360
rect 263048 325712 263100 325718
rect 263048 325654 263100 325660
rect 264256 316034 264284 329990
rect 264900 329882 264928 329990
rect 264900 329854 265020 329882
rect 264992 326466 265020 329854
rect 264980 326460 265032 326466
rect 264980 326402 265032 326408
rect 263888 316006 264284 316034
rect 262956 311228 263008 311234
rect 262956 311170 263008 311176
rect 263888 309874 263916 316006
rect 263876 309868 263928 309874
rect 263876 309810 263928 309816
rect 265084 308514 265112 329990
rect 265452 327944 265480 329990
rect 265176 327916 265480 327944
rect 265176 323610 265204 327916
rect 265912 327842 265940 329990
rect 265452 327814 265940 327842
rect 265164 323604 265216 323610
rect 265164 323546 265216 323552
rect 265072 308508 265124 308514
rect 265072 308450 265124 308456
rect 263508 95940 263560 95946
rect 263508 95882 263560 95888
rect 263520 6914 263548 95882
rect 265452 13122 265480 327814
rect 266372 327690 266400 329990
rect 266740 327842 266768 329990
rect 266464 327814 266768 327842
rect 266360 327684 266412 327690
rect 266360 327626 266412 327632
rect 265624 327140 265676 327146
rect 265624 327082 265676 327088
rect 265440 13116 265492 13122
rect 265440 13058 265492 13064
rect 265636 7682 265664 327082
rect 266464 89010 266492 327814
rect 267108 316034 267136 329990
rect 267752 327146 267780 329990
rect 267936 327962 267964 329990
rect 268304 327978 268332 329990
rect 267924 327956 267976 327962
rect 267924 327898 267976 327904
rect 268212 327950 268332 327978
rect 267740 327140 267792 327146
rect 267740 327082 267792 327088
rect 268212 316034 268240 327950
rect 268764 327842 268792 329990
rect 266740 316006 267136 316034
rect 267936 316006 268240 316034
rect 268304 327814 268792 327842
rect 268936 327820 268988 327826
rect 266452 89004 266504 89010
rect 266452 88946 266504 88952
rect 265624 7676 265676 7682
rect 265624 7618 265676 7624
rect 263428 6886 263548 6914
rect 265808 6928 265860 6934
rect 262864 6180 262916 6186
rect 262864 6122 262916 6128
rect 263428 480 263456 6886
rect 265808 6870 265860 6876
rect 265820 480 265848 6870
rect 266740 4894 266768 316006
rect 267936 6254 267964 316006
rect 268304 26994 268332 327814
rect 268936 327762 268988 327768
rect 268948 327146 268976 327762
rect 269132 327350 269160 329990
rect 269500 327842 269528 329990
rect 269224 327814 269528 327842
rect 269120 327344 269172 327350
rect 269120 327286 269172 327292
rect 268384 327140 268436 327146
rect 268384 327082 268436 327088
rect 268936 327140 268988 327146
rect 268936 327082 268988 327088
rect 268396 294642 268424 327082
rect 268384 294636 268436 294642
rect 268384 294578 268436 294584
rect 268292 26988 268344 26994
rect 268292 26930 268344 26936
rect 269224 8362 269252 327814
rect 269960 316034 269988 329990
rect 270512 327842 270540 329990
rect 269500 316006 269988 316034
rect 270420 327814 270540 327842
rect 269212 8356 269264 8362
rect 269212 8298 269264 8304
rect 269500 6934 269528 316006
rect 269488 6928 269540 6934
rect 269488 6870 269540 6876
rect 267924 6248 267976 6254
rect 267924 6190 267976 6196
rect 266728 4888 266780 4894
rect 266728 4830 266780 4836
rect 270420 3534 270448 327814
rect 271340 327690 271368 330126
rect 271328 327684 271380 327690
rect 271328 327626 271380 327632
rect 271708 9654 271736 330126
rect 272076 327962 272104 330126
rect 272536 328098 272564 330126
rect 272524 328092 272576 328098
rect 272524 328034 272576 328040
rect 272064 327956 272116 327962
rect 272064 327898 272116 327904
rect 272904 327894 272932 330126
rect 272996 329990 273102 330018
rect 272892 327888 272944 327894
rect 272892 327830 272944 327836
rect 271788 327684 271840 327690
rect 271788 327626 271840 327632
rect 271696 9648 271748 9654
rect 271696 9590 271748 9596
rect 271800 4214 271828 327626
rect 272996 11830 273024 329990
rect 273168 327956 273220 327962
rect 273168 327898 273220 327904
rect 273076 327888 273128 327894
rect 273076 327830 273128 327836
rect 272984 11824 273036 11830
rect 272984 11766 273036 11772
rect 273088 7682 273116 327830
rect 273076 7676 273128 7682
rect 273076 7618 273128 7624
rect 273180 4894 273208 327898
rect 273732 327554 273760 330126
rect 274100 327690 274128 330126
rect 274088 327684 274140 327690
rect 274088 327626 274140 327632
rect 273720 327548 273772 327554
rect 273720 327490 273772 327496
rect 274376 17270 274404 330126
rect 274548 327684 274600 327690
rect 274548 327626 274600 327632
rect 274456 327548 274508 327554
rect 274456 327490 274508 327496
rect 274364 17264 274416 17270
rect 274364 17206 274416 17212
rect 274468 13122 274496 327490
rect 274456 13116 274508 13122
rect 274456 13058 274508 13064
rect 274560 8974 274588 327626
rect 274928 326398 274956 330126
rect 275020 329990 275126 330018
rect 274916 326392 274968 326398
rect 274916 326334 274968 326340
rect 275020 324970 275048 329990
rect 275008 324964 275060 324970
rect 275008 324906 275060 324912
rect 275756 14482 275784 330126
rect 275848 329990 275954 330018
rect 275848 15910 275876 329990
rect 276584 327418 276612 330126
rect 276952 327962 276980 330126
rect 276940 327956 276992 327962
rect 276940 327898 276992 327904
rect 276664 327820 276716 327826
rect 276664 327762 276716 327768
rect 276572 327412 276624 327418
rect 276572 327354 276624 327360
rect 276676 18630 276704 327762
rect 277228 251870 277256 330126
rect 277504 329990 277610 330018
rect 277688 329990 277978 330018
rect 278056 329990 278438 330018
rect 277400 328024 277452 328030
rect 277400 327966 277452 327972
rect 277308 327412 277360 327418
rect 277308 327354 277360 327360
rect 277216 251864 277268 251870
rect 277216 251806 277268 251812
rect 277320 18630 277348 327354
rect 277412 320958 277440 327966
rect 277504 323678 277532 329990
rect 277688 328030 277716 329990
rect 277676 328024 277728 328030
rect 277676 327966 277728 327972
rect 277492 323672 277544 323678
rect 277492 323614 277544 323620
rect 277400 320952 277452 320958
rect 277400 320894 277452 320900
rect 278056 319530 278084 329990
rect 278976 327690 279004 330126
rect 278964 327684 279016 327690
rect 278964 327626 279016 327632
rect 279436 327554 279464 330126
rect 279516 328024 279568 328030
rect 279516 327966 279568 327972
rect 279424 327548 279476 327554
rect 279424 327490 279476 327496
rect 279424 327344 279476 327350
rect 279424 327286 279476 327292
rect 278044 319524 278096 319530
rect 278044 319466 278096 319472
rect 279436 19990 279464 327286
rect 279528 28286 279556 327966
rect 279804 327894 279832 330126
rect 279896 329990 280002 330018
rect 279792 327888 279844 327894
rect 279792 327830 279844 327836
rect 279896 327842 279924 329990
rect 280068 327888 280120 327894
rect 279896 327814 280016 327842
rect 280068 327830 280120 327836
rect 279792 327684 279844 327690
rect 279792 327626 279844 327632
rect 279804 318170 279832 327626
rect 279884 327548 279936 327554
rect 279884 327490 279936 327496
rect 279792 318164 279844 318170
rect 279792 318106 279844 318112
rect 279896 316810 279924 327490
rect 279884 316804 279936 316810
rect 279884 316746 279936 316752
rect 279988 315314 280016 327814
rect 279976 315308 280028 315314
rect 279976 315250 280028 315256
rect 280080 217326 280108 327830
rect 280632 327418 280660 330126
rect 280804 328092 280856 328098
rect 280804 328034 280856 328040
rect 280620 327412 280672 327418
rect 280620 327354 280672 327360
rect 280068 217320 280120 217326
rect 280068 217262 280120 217268
rect 279516 28280 279568 28286
rect 279516 28222 279568 28228
rect 279424 19984 279476 19990
rect 279424 19926 279476 19932
rect 276664 18624 276716 18630
rect 276664 18566 276716 18572
rect 277308 18624 277360 18630
rect 277308 18566 277360 18572
rect 275836 15904 275888 15910
rect 275836 15846 275888 15852
rect 275744 14476 275796 14482
rect 275744 14418 275796 14424
rect 276480 9648 276532 9654
rect 276480 9590 276532 9596
rect 274548 8968 274600 8974
rect 274548 8910 274600 8916
rect 273168 4888 273220 4894
rect 273168 4830 273220 4836
rect 271788 4208 271840 4214
rect 271788 4150 271840 4156
rect 272892 4208 272944 4214
rect 272892 4150 272944 4156
rect 269304 3528 269356 3534
rect 269304 3470 269356 3476
rect 270408 3528 270460 3534
rect 270408 3470 270460 3476
rect 270500 3528 270552 3534
rect 270500 3470 270552 3476
rect 267004 3460 267056 3466
rect 267004 3402 267056 3408
rect 267016 480 267044 3402
rect 269316 480 269344 3470
rect 270512 480 270540 3470
rect 272904 480 272932 4150
rect 274088 3596 274140 3602
rect 274088 3538 274140 3544
rect 274100 480 274128 3538
rect 276492 480 276520 9590
rect 280068 4888 280120 4894
rect 280068 4830 280120 4836
rect 277676 3732 277728 3738
rect 277676 3674 277728 3680
rect 277688 480 277716 3674
rect 280080 480 280108 4830
rect 280816 4214 280844 328034
rect 281092 327842 281120 330126
rect 281092 327814 281396 327842
rect 281264 327412 281316 327418
rect 281264 327354 281316 327360
rect 281276 6254 281304 327354
rect 281264 6248 281316 6254
rect 281264 6190 281316 6196
rect 281368 6186 281396 327814
rect 281356 6180 281408 6186
rect 281356 6122 281408 6128
rect 280804 4208 280856 4214
rect 280804 4150 280856 4156
rect 281264 3800 281316 3806
rect 281264 3742 281316 3748
rect 281276 480 281304 3742
rect 281460 3670 281488 330126
rect 281552 329990 281658 330018
rect 281828 329990 282026 330018
rect 282104 329990 282486 330018
rect 282564 329990 282854 330018
rect 283116 329990 283314 330018
rect 283392 329990 283682 330018
rect 283760 329990 284050 330018
rect 284404 329990 284510 330018
rect 284588 329990 284878 330018
rect 285048 329990 285338 330018
rect 281552 327826 281580 329990
rect 281724 327888 281776 327894
rect 281724 327830 281776 327836
rect 281540 327820 281592 327826
rect 281540 327762 281592 327768
rect 281736 286346 281764 327830
rect 281828 327758 281856 329990
rect 281816 327752 281868 327758
rect 281816 327694 281868 327700
rect 282104 287706 282132 329990
rect 282564 327894 282592 329990
rect 282552 327888 282604 327894
rect 282552 327830 282604 327836
rect 283012 327888 283064 327894
rect 283012 327830 283064 327836
rect 282920 327820 282972 327826
rect 282920 327762 282972 327768
rect 282092 287700 282144 287706
rect 282092 287642 282144 287648
rect 281724 286340 281776 286346
rect 281724 286282 281776 286288
rect 282932 37942 282960 327762
rect 283024 283626 283052 327830
rect 283116 284986 283144 329990
rect 283392 327894 283420 329990
rect 283380 327888 283432 327894
rect 283380 327830 283432 327836
rect 283760 327826 283788 329990
rect 283748 327820 283800 327826
rect 283748 327762 283800 327768
rect 284404 325694 284432 329990
rect 284404 325666 284524 325694
rect 283104 284980 283156 284986
rect 283104 284922 283156 284928
rect 283012 283620 283064 283626
rect 283012 283562 283064 283568
rect 282920 37936 282972 37942
rect 282920 37878 282972 37884
rect 284496 10334 284524 325666
rect 284588 42090 284616 329990
rect 284944 327888 284996 327894
rect 284944 327830 284996 327836
rect 284956 300150 284984 327830
rect 285048 327350 285076 329990
rect 285784 327894 285812 330126
rect 285876 329990 286166 330018
rect 286244 329990 286534 330018
rect 286612 329990 286902 330018
rect 287164 329990 287362 330018
rect 287440 329990 287730 330018
rect 287808 329990 288190 330018
rect 288452 329990 288558 330018
rect 288636 329990 288926 330018
rect 289096 329990 289386 330018
rect 289464 329990 289754 330018
rect 289832 329990 290214 330018
rect 290292 329990 290582 330018
rect 290752 329990 291042 330018
rect 291212 329990 291410 330018
rect 291488 329990 291778 330018
rect 291856 329990 292238 330018
rect 285876 328166 285904 329990
rect 285864 328160 285916 328166
rect 285864 328102 285916 328108
rect 285772 327888 285824 327894
rect 285772 327830 285824 327836
rect 285772 327752 285824 327758
rect 285772 327694 285824 327700
rect 285036 327344 285088 327350
rect 285036 327286 285088 327292
rect 284944 300144 284996 300150
rect 284944 300086 284996 300092
rect 285784 298790 285812 327694
rect 286244 316034 286272 329990
rect 286612 327758 286640 329990
rect 286600 327752 286652 327758
rect 286600 327694 286652 327700
rect 287164 327146 287192 329990
rect 286324 327140 286376 327146
rect 286324 327082 286376 327088
rect 287152 327140 287204 327146
rect 287152 327082 287204 327088
rect 285876 316006 286272 316034
rect 285772 298784 285824 298790
rect 285772 298726 285824 298732
rect 284576 42084 284628 42090
rect 284576 42026 284628 42032
rect 285876 21418 285904 316006
rect 286336 22778 286364 327082
rect 287440 326482 287468 329990
rect 287808 327978 287836 329990
rect 287164 326454 287468 326482
rect 287624 327950 287836 327978
rect 287164 25566 287192 326454
rect 287624 316034 287652 327950
rect 288452 327894 288480 329990
rect 287796 327888 287848 327894
rect 287796 327830 287848 327836
rect 288440 327888 288492 327894
rect 288440 327830 288492 327836
rect 287704 327684 287756 327690
rect 287704 327626 287756 327632
rect 287440 316006 287652 316034
rect 287152 25560 287204 25566
rect 287152 25502 287204 25508
rect 287440 24138 287468 316006
rect 287716 296002 287744 327626
rect 287808 297430 287836 327830
rect 288636 327690 288664 329990
rect 289096 328030 289124 329990
rect 289084 328024 289136 328030
rect 289084 327966 289136 327972
rect 288624 327684 288676 327690
rect 288624 327626 288676 327632
rect 289464 316034 289492 329990
rect 288636 316006 289492 316034
rect 287796 297424 287848 297430
rect 287796 297366 287848 297372
rect 287704 295996 287756 296002
rect 287704 295938 287756 295944
rect 288636 293282 288664 316006
rect 288624 293276 288676 293282
rect 288624 293218 288676 293224
rect 289832 32434 289860 329990
rect 289912 327820 289964 327826
rect 289912 327762 289964 327768
rect 289924 290494 289952 327762
rect 290292 316034 290320 329990
rect 290464 327888 290516 327894
rect 290464 327830 290516 327836
rect 290016 316006 290320 316034
rect 290016 291854 290044 316006
rect 290004 291848 290056 291854
rect 290004 291790 290056 291796
rect 289912 290488 289964 290494
rect 289912 290430 289964 290436
rect 289820 32428 289872 32434
rect 289820 32370 289872 32376
rect 290476 31074 290504 327830
rect 290752 327826 290780 329990
rect 291212 327894 291240 329990
rect 291200 327888 291252 327894
rect 291200 327830 291252 327836
rect 290740 327820 290792 327826
rect 290740 327762 290792 327768
rect 291488 33794 291516 329990
rect 291856 327842 291884 329990
rect 292684 327894 292712 330126
rect 292776 329990 293066 330018
rect 293144 329990 293434 330018
rect 293512 329990 293802 330018
rect 294064 329990 294262 330018
rect 294340 329990 294630 330018
rect 294708 329990 295090 330018
rect 295352 329990 295458 330018
rect 295628 329990 295918 330018
rect 295996 329990 296286 330018
rect 296364 329990 296654 330018
rect 296732 329990 297114 330018
rect 297192 329990 297482 330018
rect 297560 329990 297942 330018
rect 298204 329990 298310 330018
rect 298388 329990 298678 330018
rect 298756 329990 299138 330018
rect 291580 327814 291884 327842
rect 291936 327888 291988 327894
rect 291936 327830 291988 327836
rect 292672 327888 292724 327894
rect 292672 327830 292724 327836
rect 291580 35222 291608 327814
rect 291844 327616 291896 327622
rect 291844 327558 291896 327564
rect 291568 35216 291620 35222
rect 291568 35158 291620 35164
rect 291476 33788 291528 33794
rect 291476 33730 291528 33736
rect 290464 31068 290516 31074
rect 290464 31010 290516 31016
rect 287428 24132 287480 24138
rect 287428 24074 287480 24080
rect 286324 22772 286376 22778
rect 286324 22714 286376 22720
rect 285864 21412 285916 21418
rect 285864 21354 285916 21360
rect 290740 11824 290792 11830
rect 290740 11766 290792 11772
rect 284484 10328 284536 10334
rect 284484 10270 284536 10276
rect 287152 7676 287204 7682
rect 287152 7618 287204 7624
rect 283656 4208 283708 4214
rect 283656 4150 283708 4156
rect 281448 3664 281500 3670
rect 281448 3606 281500 3612
rect 283668 480 283696 4150
rect 284760 3868 284812 3874
rect 284760 3810 284812 3816
rect 284772 480 284800 3810
rect 287164 480 287192 7618
rect 288348 3936 288400 3942
rect 288348 3878 288400 3884
rect 288360 480 288388 3878
rect 290752 480 290780 11766
rect 291856 7614 291884 327558
rect 291948 289202 291976 327830
rect 292672 327752 292724 327758
rect 292672 327694 292724 327700
rect 291936 289196 291988 289202
rect 291936 289138 291988 289144
rect 292684 39370 292712 327694
rect 292776 322318 292804 329990
rect 293144 327758 293172 329990
rect 293132 327752 293184 327758
rect 293132 327694 293184 327700
rect 292764 322312 292816 322318
rect 292764 322254 292816 322260
rect 293512 316034 293540 329990
rect 293960 328024 294012 328030
rect 293960 327966 294012 327972
rect 292868 316006 293540 316034
rect 292672 39364 292724 39370
rect 292672 39306 292724 39312
rect 292868 36582 292896 316006
rect 292856 36576 292908 36582
rect 292856 36518 292908 36524
rect 291844 7608 291896 7614
rect 291844 7550 291896 7556
rect 293972 4826 294000 327966
rect 294064 11762 294092 329990
rect 294340 328030 294368 329990
rect 294328 328024 294380 328030
rect 294328 327966 294380 327972
rect 294708 327842 294736 329990
rect 294340 327814 294736 327842
rect 294340 29714 294368 327814
rect 294604 327684 294656 327690
rect 294604 327626 294656 327632
rect 294616 304298 294644 327626
rect 295352 327622 295380 329990
rect 295524 327888 295576 327894
rect 295524 327830 295576 327836
rect 295340 327616 295392 327622
rect 295340 327558 295392 327564
rect 294604 304292 294656 304298
rect 294604 304234 294656 304240
rect 295536 95946 295564 327830
rect 295628 327690 295656 329990
rect 295616 327684 295668 327690
rect 295616 327626 295668 327632
rect 295996 316034 296024 329990
rect 296364 327894 296392 329990
rect 296352 327888 296404 327894
rect 296352 327830 296404 327836
rect 295720 316006 296024 316034
rect 295720 312594 295748 316006
rect 295708 312588 295760 312594
rect 295708 312530 295760 312536
rect 295524 95940 295576 95946
rect 295524 95882 295576 95888
rect 294328 29708 294380 29714
rect 294328 29650 294380 29656
rect 294328 13116 294380 13122
rect 294328 13058 294380 13064
rect 294052 11756 294104 11762
rect 294052 11698 294104 11704
rect 293960 4820 294012 4826
rect 293960 4762 294012 4768
rect 291936 4004 291988 4010
rect 291936 3946 291988 3952
rect 291948 480 291976 3946
rect 294340 480 294368 13058
rect 295524 4072 295576 4078
rect 295524 4014 295576 4020
rect 295536 480 295564 4014
rect 296732 3466 296760 329990
rect 297192 327842 297220 329990
rect 296824 327814 297220 327842
rect 296824 3534 296852 327814
rect 297560 316034 297588 329990
rect 298100 327888 298152 327894
rect 298100 327830 298152 327836
rect 296916 316006 297588 316034
rect 296916 3602 296944 316006
rect 297916 8968 297968 8974
rect 297916 8910 297968 8916
rect 296904 3596 296956 3602
rect 296904 3538 296956 3544
rect 296812 3528 296864 3534
rect 296812 3470 296864 3476
rect 296720 3460 296772 3466
rect 296720 3402 296772 3408
rect 297928 480 297956 8910
rect 298112 3806 298140 327830
rect 298100 3800 298152 3806
rect 298100 3742 298152 3748
rect 298204 3738 298232 329990
rect 298388 327894 298416 329990
rect 298376 327888 298428 327894
rect 298376 327830 298428 327836
rect 298756 316034 298784 329990
rect 299584 327842 299612 330126
rect 298388 316006 298784 316034
rect 299492 327814 299612 327842
rect 299676 329990 299966 330018
rect 300044 329990 300334 330018
rect 300412 329990 300794 330018
rect 298388 3874 298416 316006
rect 299492 3942 299520 327814
rect 299572 327752 299624 327758
rect 299572 327694 299624 327700
rect 299584 4078 299612 327694
rect 299572 4072 299624 4078
rect 299572 4014 299624 4020
rect 299676 4010 299704 329990
rect 300044 327758 300072 329990
rect 300032 327752 300084 327758
rect 300032 327694 300084 327700
rect 300412 316034 300440 329990
rect 300952 328024 301004 328030
rect 300952 327966 301004 327972
rect 300964 322250 300992 327966
rect 301332 327554 301360 330126
rect 301792 327842 301820 330126
rect 301884 329990 301990 330018
rect 301884 328030 301912 329990
rect 302620 328166 302648 330126
rect 302608 328160 302660 328166
rect 302608 328102 302660 328108
rect 301872 328024 301924 328030
rect 301872 327966 301924 327972
rect 301792 327814 302188 327842
rect 301320 327548 301372 327554
rect 301320 327490 301372 327496
rect 302056 327548 302108 327554
rect 302056 327490 302108 327496
rect 300952 322244 301004 322250
rect 300952 322186 301004 322192
rect 299768 316006 300440 316034
rect 299664 4004 299716 4010
rect 299664 3946 299716 3952
rect 299480 3936 299532 3942
rect 299480 3878 299532 3884
rect 298376 3868 298428 3874
rect 298376 3810 298428 3816
rect 298192 3732 298244 3738
rect 298192 3674 298244 3680
rect 299768 3534 299796 316006
rect 300860 17264 300912 17270
rect 300860 17206 300912 17212
rect 300872 16574 300900 17206
rect 300872 16546 301452 16574
rect 299112 3528 299164 3534
rect 299112 3470 299164 3476
rect 299756 3528 299808 3534
rect 299756 3470 299808 3476
rect 299124 480 299152 3470
rect 301424 480 301452 16546
rect 302068 3534 302096 327490
rect 302056 3528 302108 3534
rect 302056 3470 302108 3476
rect 302160 3194 302188 327814
rect 302988 327758 303016 330126
rect 302976 327752 303028 327758
rect 302976 327694 303028 327700
rect 302608 3528 302660 3534
rect 302608 3470 302660 3476
rect 302148 3188 302200 3194
rect 302148 3130 302200 3136
rect 302620 480 302648 3470
rect 303356 3398 303384 330126
rect 303448 329990 303554 330018
rect 303448 327842 303476 329990
rect 303448 327814 303568 327842
rect 303436 327752 303488 327758
rect 303436 327694 303488 327700
rect 303448 3466 303476 327694
rect 303540 3942 303568 327814
rect 304184 327622 304212 330126
rect 304172 327616 304224 327622
rect 304172 327558 304224 327564
rect 304644 327554 304672 330126
rect 304736 329990 304842 330018
rect 304632 327548 304684 327554
rect 304632 327490 304684 327496
rect 303528 3936 303580 3942
rect 303528 3878 303580 3884
rect 304736 3738 304764 329990
rect 304816 327616 304868 327622
rect 304816 327558 304868 327564
rect 304828 4078 304856 327558
rect 304908 327548 304960 327554
rect 304908 327490 304960 327496
rect 304816 4072 304868 4078
rect 304816 4014 304868 4020
rect 304920 4010 304948 327490
rect 305472 327418 305500 330126
rect 305460 327412 305512 327418
rect 305460 327354 305512 327360
rect 305092 326392 305144 326398
rect 305092 326334 305144 326340
rect 305104 6914 305132 326334
rect 305840 325694 305868 330126
rect 306208 328030 306236 330126
rect 306196 328024 306248 328030
rect 306196 327966 306248 327972
rect 306668 327418 306696 330126
rect 307036 328098 307064 330126
rect 307024 328092 307076 328098
rect 307024 328034 307076 328040
rect 307496 327826 307524 330126
rect 307588 329990 307694 330018
rect 307588 327842 307616 329990
rect 307484 327820 307536 327826
rect 307588 327814 307708 327842
rect 307484 327762 307536 327768
rect 306288 327412 306340 327418
rect 306288 327354 306340 327360
rect 306656 327412 306708 327418
rect 306656 327354 306708 327360
rect 307576 327412 307628 327418
rect 307576 327354 307628 327360
rect 305840 325666 306236 325694
rect 305012 6886 305132 6914
rect 304908 4004 304960 4010
rect 304908 3946 304960 3952
rect 304724 3732 304776 3738
rect 304724 3674 304776 3680
rect 303436 3460 303488 3466
rect 303436 3402 303488 3408
rect 303344 3392 303396 3398
rect 303344 3334 303396 3340
rect 305012 480 305040 6886
rect 306208 3806 306236 325666
rect 306300 3874 306328 327354
rect 306288 3868 306340 3874
rect 306288 3810 306340 3816
rect 306196 3800 306248 3806
rect 306196 3742 306248 3748
rect 307588 3602 307616 327354
rect 307576 3596 307628 3602
rect 307576 3538 307628 3544
rect 307680 3330 307708 327814
rect 308232 327758 308260 330126
rect 308220 327752 308272 327758
rect 308220 327694 308272 327700
rect 308692 327554 308720 330126
rect 308680 327548 308732 327554
rect 308680 327490 308732 327496
rect 307760 324964 307812 324970
rect 307760 324906 307812 324912
rect 307772 16574 307800 324906
rect 307772 16546 308628 16574
rect 307668 3324 307720 3330
rect 307668 3266 307720 3272
rect 306196 3188 306248 3194
rect 306196 3130 306248 3136
rect 306208 480 306236 3130
rect 308600 480 308628 16546
rect 308968 4826 308996 330126
rect 309048 327548 309100 327554
rect 309048 327490 309100 327496
rect 308956 4820 309008 4826
rect 308956 4762 309008 4768
rect 309060 3534 309088 327490
rect 309336 326398 309364 330126
rect 309428 329990 309718 330018
rect 309324 326392 309376 326398
rect 309324 326334 309376 326340
rect 309428 324970 309456 329990
rect 309416 324964 309468 324970
rect 309416 324906 309468 324912
rect 309140 322244 309192 322250
rect 309140 322186 309192 322192
rect 309152 16574 309180 322186
rect 309152 16546 309824 16574
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309796 480 309824 16546
rect 310256 7614 310284 330126
rect 310624 323610 310652 330126
rect 311084 327418 311112 330126
rect 311452 327554 311480 330126
rect 311544 329990 311742 330018
rect 311440 327548 311492 327554
rect 311440 327490 311492 327496
rect 311072 327412 311124 327418
rect 311072 327354 311124 327360
rect 310612 323604 310664 323610
rect 310612 323546 310664 323552
rect 311544 309806 311572 329990
rect 312372 328234 312400 330126
rect 312360 328228 312412 328234
rect 312360 328170 312412 328176
rect 312544 328160 312596 328166
rect 312544 328102 312596 328108
rect 311716 327548 311768 327554
rect 311716 327490 311768 327496
rect 311624 327412 311676 327418
rect 311624 327354 311676 327360
rect 311636 313954 311664 327354
rect 311624 313948 311676 313954
rect 311624 313890 311676 313896
rect 311728 312594 311756 327490
rect 311716 312588 311768 312594
rect 311716 312530 311768 312536
rect 311532 309800 311584 309806
rect 311532 309742 311584 309748
rect 312176 14476 312228 14482
rect 312176 14418 312228 14424
rect 310244 7608 310296 7614
rect 310244 7550 310296 7556
rect 312188 480 312216 14418
rect 312556 4214 312584 328102
rect 312740 325694 312768 330126
rect 313108 327842 313136 330126
rect 313108 327814 313228 327842
rect 312740 325666 313136 325694
rect 313108 308446 313136 325666
rect 313096 308440 313148 308446
rect 313096 308382 313148 308388
rect 313200 14482 313228 327814
rect 313384 320890 313412 330126
rect 313568 329990 313766 330018
rect 313372 320884 313424 320890
rect 313372 320826 313424 320832
rect 313568 319462 313596 329990
rect 314396 328370 314424 330126
rect 314488 329990 314594 330018
rect 314384 328364 314436 328370
rect 314384 328306 314436 328312
rect 314488 325694 314516 329990
rect 315224 327894 315252 330126
rect 315212 327888 315264 327894
rect 315212 327830 315264 327836
rect 315592 327486 315620 330126
rect 315764 327888 315816 327894
rect 315764 327830 315816 327836
rect 315580 327480 315632 327486
rect 315580 327422 315632 327428
rect 314488 325666 314608 325694
rect 313556 319456 313608 319462
rect 313556 319398 313608 319404
rect 314580 307086 314608 325666
rect 314568 307080 314620 307086
rect 314568 307022 314620 307028
rect 315776 305658 315804 327830
rect 315764 305652 315816 305658
rect 315764 305594 315816 305600
rect 315868 304298 315896 330126
rect 316420 327690 316448 330126
rect 316408 327684 316460 327690
rect 316408 327626 316460 327632
rect 316788 327554 316816 330126
rect 317144 327684 317196 327690
rect 317144 327626 317196 327632
rect 316776 327548 316828 327554
rect 316776 327490 316828 327496
rect 315948 327480 316000 327486
rect 315948 327422 316000 327428
rect 315856 304292 315908 304298
rect 315856 304234 315908 304240
rect 315960 15910 315988 327422
rect 317156 302938 317184 327626
rect 317144 302932 317196 302938
rect 317144 302874 317196 302880
rect 317248 301510 317276 330126
rect 317616 327962 317644 330126
rect 317604 327956 317656 327962
rect 317604 327898 317656 327904
rect 317984 327690 318012 330126
rect 318444 328114 318472 330126
rect 318444 328086 318656 328114
rect 318432 327956 318484 327962
rect 318432 327898 318484 327904
rect 317972 327684 318024 327690
rect 317972 327626 318024 327632
rect 317328 327548 317380 327554
rect 317328 327490 317380 327496
rect 317236 301504 317288 301510
rect 317236 301446 317288 301452
rect 317340 133210 317368 327490
rect 318444 318102 318472 327898
rect 318524 327684 318576 327690
rect 318524 327626 318576 327632
rect 318432 318096 318484 318102
rect 318432 318038 318484 318044
rect 318536 316742 318564 327626
rect 318524 316736 318576 316742
rect 318524 316678 318576 316684
rect 318628 300150 318656 328086
rect 318616 300144 318668 300150
rect 318616 300086 318668 300092
rect 318720 298790 318748 330126
rect 319272 327690 319300 330126
rect 319640 327842 319668 330126
rect 319640 327814 320036 327842
rect 319260 327684 319312 327690
rect 319260 327626 319312 327632
rect 319904 327684 319956 327690
rect 319904 327626 319956 327632
rect 318708 298784 318760 298790
rect 318708 298726 318760 298732
rect 319916 297430 319944 327626
rect 319904 297424 319956 297430
rect 319904 297366 319956 297372
rect 320008 296002 320036 327814
rect 319996 295996 320048 296002
rect 319996 295938 320048 295944
rect 317328 133204 317380 133210
rect 317328 133146 317380 133152
rect 318800 18624 318852 18630
rect 318800 18566 318852 18572
rect 318812 16574 318840 18566
rect 318812 16546 319300 16574
rect 315764 15904 315816 15910
rect 315764 15846 315816 15852
rect 315948 15904 316000 15910
rect 315948 15846 316000 15852
rect 313188 14476 313240 14482
rect 313188 14418 313240 14424
rect 312544 4208 312596 4214
rect 312544 4150 312596 4156
rect 313372 4208 313424 4214
rect 313372 4150 313424 4156
rect 313384 480 313412 4150
rect 315776 480 315804 15846
rect 316960 3460 317012 3466
rect 316960 3402 317012 3408
rect 316972 480 317000 3402
rect 319272 480 319300 16546
rect 320100 3466 320128 330126
rect 320916 328364 320968 328370
rect 320916 328306 320968 328312
rect 320824 327616 320876 327622
rect 320824 327558 320876 327564
rect 320836 9654 320864 327558
rect 320928 10334 320956 328306
rect 322216 41410 322244 336767
rect 322308 77246 322336 339374
rect 322400 135250 322428 352543
rect 322492 171086 322520 357983
rect 322584 229090 322612 366143
rect 322676 264926 322704 368863
rect 322768 322930 322796 398919
rect 334624 396092 334676 396098
rect 334624 396034 334676 396040
rect 333244 360256 333296 360262
rect 333244 360198 333296 360204
rect 326344 355156 326396 355162
rect 326344 355098 326396 355104
rect 323584 328228 323636 328234
rect 323584 328170 323636 328176
rect 322756 322924 322808 322930
rect 322756 322866 322808 322872
rect 322664 264920 322716 264926
rect 322664 264862 322716 264868
rect 322572 229084 322624 229090
rect 322572 229026 322624 229032
rect 322480 171080 322532 171086
rect 322480 171022 322532 171028
rect 322388 135244 322440 135250
rect 322388 135186 322440 135192
rect 322296 77240 322348 77246
rect 322296 77182 322348 77188
rect 322204 41404 322256 41410
rect 322204 41346 322256 41352
rect 320916 10328 320968 10334
rect 320916 10270 320968 10276
rect 320824 9648 320876 9654
rect 320824 9590 320876 9596
rect 322848 9648 322900 9654
rect 322848 9590 322900 9596
rect 320088 3460 320140 3466
rect 320088 3402 320140 3408
rect 320456 3392 320508 3398
rect 320456 3334 320508 3340
rect 320468 480 320496 3334
rect 322860 480 322888 9590
rect 323596 8974 323624 328170
rect 326356 252550 326384 355098
rect 327724 345092 327776 345098
rect 327724 345034 327776 345040
rect 326344 252544 326396 252550
rect 326344 252486 326396 252492
rect 325700 251864 325752 251870
rect 325700 251806 325752 251812
rect 325712 16574 325740 251806
rect 327736 88330 327764 345034
rect 329840 323672 329892 323678
rect 329840 323614 329892 323620
rect 327724 88324 327776 88330
rect 327724 88266 327776 88272
rect 329852 16574 329880 323614
rect 332600 320952 332652 320958
rect 332600 320894 332652 320900
rect 332612 16574 332640 320894
rect 333256 182170 333284 360198
rect 334636 276010 334664 396034
rect 388456 383654 388484 498170
rect 391216 386374 391244 545090
rect 393976 416770 394004 603094
rect 395344 462392 395396 462398
rect 395344 462334 395396 462340
rect 393964 416764 394016 416770
rect 393964 416706 394016 416712
rect 394056 415472 394108 415478
rect 394056 415414 394108 415420
rect 394068 405686 394096 415414
rect 395356 408474 395384 462334
rect 397472 423230 397500 703520
rect 413664 700398 413692 703520
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 462332 700330 462360 703520
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 478524 683114 478552 703520
rect 477512 683086 478552 683114
rect 397460 423224 397512 423230
rect 397460 423166 397512 423172
rect 477512 423162 477540 683086
rect 477500 423156 477552 423162
rect 477500 423098 477552 423104
rect 527192 423026 527220 703520
rect 543476 683114 543504 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 686352 580318 686361
rect 580262 686287 580318 686296
rect 542372 683086 543504 683114
rect 527180 423020 527232 423026
rect 527180 422962 527232 422968
rect 542372 422958 542400 683086
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 579802 557288 579858 557297
rect 579802 557223 579858 557232
rect 579816 556238 579844 557223
rect 579804 556232 579856 556238
rect 579804 556174 579856 556180
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 579802 510368 579858 510377
rect 579802 510303 579858 510312
rect 579816 509318 579844 510303
rect 579804 509312 579856 509318
rect 579804 509254 579856 509260
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 579802 463448 579858 463457
rect 579802 463383 579858 463392
rect 579816 462398 579844 463383
rect 579804 462392 579856 462398
rect 579804 462334 579856 462340
rect 542360 422952 542412 422958
rect 542360 422894 542412 422900
rect 579618 416528 579674 416537
rect 579618 416463 579674 416472
rect 579632 415478 579660 416463
rect 579620 415472 579672 415478
rect 579620 415414 579672 415420
rect 395344 408468 395396 408474
rect 395344 408410 395396 408416
rect 394056 405680 394108 405686
rect 394056 405622 394108 405628
rect 580276 394670 580304 686287
rect 580354 639432 580410 639441
rect 580354 639367 580410 639376
rect 580264 394664 580316 394670
rect 580264 394606 580316 394612
rect 580368 391950 580396 639367
rect 580446 592512 580502 592521
rect 580446 592447 580502 592456
rect 580356 391944 580408 391950
rect 580356 391886 580408 391892
rect 580460 389162 580488 592447
rect 580538 451752 580594 451761
rect 580538 451687 580594 451696
rect 580448 389156 580500 389162
rect 580448 389098 580500 389104
rect 391204 386368 391256 386374
rect 391204 386310 391256 386316
rect 388444 383648 388496 383654
rect 388444 383590 388496 383596
rect 580552 380866 580580 451687
rect 580630 404832 580686 404841
rect 580630 404767 580686 404776
rect 580540 380860 580592 380866
rect 580540 380802 580592 380808
rect 580644 378146 580672 404767
rect 580632 378140 580684 378146
rect 580632 378082 580684 378088
rect 355324 371272 355376 371278
rect 355324 371214 355376 371220
rect 348424 362976 348476 362982
rect 348424 362918 348476 362924
rect 341524 349172 341576 349178
rect 341524 349114 341576 349120
rect 340144 334008 340196 334014
rect 340144 333950 340196 333956
rect 336740 319524 336792 319530
rect 336740 319466 336792 319472
rect 334624 276004 334676 276010
rect 334624 275946 334676 275952
rect 333244 182164 333296 182170
rect 333244 182106 333296 182112
rect 336752 16574 336780 319466
rect 339500 318164 339552 318170
rect 339500 318106 339552 318112
rect 325712 16546 326476 16574
rect 329852 16546 330064 16574
rect 332612 16546 333652 16574
rect 336752 16546 337148 16574
rect 323584 8968 323636 8974
rect 323584 8910 323636 8916
rect 324044 4140 324096 4146
rect 324044 4082 324096 4088
rect 324056 480 324084 4082
rect 326448 480 326476 16546
rect 327632 4072 327684 4078
rect 327632 4014 327684 4020
rect 327644 480 327672 4014
rect 330036 480 330064 16546
rect 331220 4004 331272 4010
rect 331220 3946 331272 3952
rect 331232 480 331260 3946
rect 333624 480 333652 16546
rect 334716 3936 334768 3942
rect 334716 3878 334768 3884
rect 334728 480 334756 3878
rect 337120 480 337148 16546
rect 338304 3868 338356 3874
rect 338304 3810 338356 3816
rect 338316 480 338344 3810
rect 339512 3398 339540 318106
rect 340156 30326 340184 333950
rect 341536 124166 341564 349114
rect 345020 328024 345072 328030
rect 345020 327966 345072 327972
rect 343640 316804 343692 316810
rect 343640 316746 343692 316752
rect 341524 124160 341576 124166
rect 341524 124102 341576 124108
rect 340144 30320 340196 30326
rect 340144 30262 340196 30268
rect 343652 16574 343680 316746
rect 345032 16574 345060 327966
rect 348436 218006 348464 362918
rect 351920 327888 351972 327894
rect 351920 327830 351972 327836
rect 350540 315308 350592 315314
rect 350540 315250 350592 315256
rect 348424 218000 348476 218006
rect 348424 217942 348476 217948
rect 347872 217320 347924 217326
rect 347872 217262 347924 217268
rect 343652 16546 344324 16574
rect 345032 16546 345520 16574
rect 341892 3800 341944 3806
rect 341892 3742 341944 3748
rect 339500 3392 339552 3398
rect 339500 3334 339552 3340
rect 340696 3392 340748 3398
rect 340696 3334 340748 3340
rect 340708 480 340736 3334
rect 341904 480 341932 3742
rect 344296 480 344324 16546
rect 345492 480 345520 16546
rect 347884 480 347912 217262
rect 350552 16574 350580 315250
rect 351932 16574 351960 327830
rect 355336 311846 355364 371214
rect 580172 369844 580224 369850
rect 580172 369786 580224 369792
rect 580184 369617 580212 369786
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 579988 358760 580040 358766
rect 579988 358702 580040 358708
rect 580000 357921 580028 358702
rect 579986 357912 580042 357921
rect 579986 357847 580042 357856
rect 384304 346452 384356 346458
rect 384304 346394 384356 346400
rect 355324 311840 355376 311846
rect 355324 311782 355376 311788
rect 384316 111790 384344 346394
rect 406384 339516 406436 339522
rect 406384 339458 406436 339464
rect 384304 111784 384356 111790
rect 384304 111726 384356 111732
rect 406396 64870 406424 339458
rect 429844 331288 429896 331294
rect 429844 331230 429896 331236
rect 406384 64864 406436 64870
rect 406384 64806 406436 64812
rect 429856 17950 429884 331230
rect 469220 327820 469272 327826
rect 469220 327762 469272 327768
rect 429844 17944 429896 17950
rect 429844 17886 429896 17892
rect 469232 16574 469260 327762
rect 477500 327752 477552 327758
rect 477500 327694 477552 327700
rect 350552 16546 351408 16574
rect 351932 16546 352604 16574
rect 469232 16546 470364 16574
rect 349068 3732 349120 3738
rect 349068 3674 349120 3680
rect 349080 480 349108 3674
rect 351380 480 351408 16546
rect 352576 480 352604 16546
rect 354956 6248 355008 6254
rect 354956 6190 355008 6196
rect 354968 480 354996 6190
rect 358544 6180 358596 6186
rect 358544 6122 358596 6128
rect 358556 480 358584 6122
rect 363328 3664 363380 3670
rect 363328 3606 363380 3612
rect 363340 480 363368 3606
rect 470336 480 470364 16546
rect 473912 3596 473964 3602
rect 473912 3538 473964 3544
rect 473924 480 473952 3538
rect 477512 480 477540 327694
rect 487160 326392 487212 326398
rect 487160 326334 487212 326340
rect 487172 16574 487200 326334
rect 491300 324964 491352 324970
rect 491300 324906 491352 324912
rect 491312 16574 491340 324906
rect 498200 323604 498252 323610
rect 498200 323546 498252 323552
rect 498212 16574 498240 323546
rect 580172 322924 580224 322930
rect 580172 322866 580224 322872
rect 580184 322697 580212 322866
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 523040 320884 523092 320890
rect 523040 320826 523092 320832
rect 502340 313948 502392 313954
rect 502340 313890 502392 313896
rect 502352 16574 502380 313890
rect 505100 312588 505152 312594
rect 505100 312530 505152 312536
rect 505112 16574 505140 312530
rect 509240 309800 509292 309806
rect 509240 309742 509292 309748
rect 509252 16574 509280 309742
rect 516140 308440 516192 308446
rect 516140 308382 516192 308388
rect 516152 16574 516180 308382
rect 523052 16574 523080 320826
rect 527180 319456 527232 319462
rect 527180 319398 527232 319404
rect 527192 16574 527220 319398
rect 558184 318096 558236 318102
rect 558184 318038 558236 318044
rect 534080 307080 534132 307086
rect 534080 307022 534132 307028
rect 534092 16574 534120 307022
rect 536840 305652 536892 305658
rect 536840 305594 536892 305600
rect 487172 16546 488212 16574
rect 491312 16546 491800 16574
rect 498212 16546 498976 16574
rect 502352 16546 502472 16574
rect 505112 16546 506060 16574
rect 509252 16546 509648 16574
rect 516152 16546 516824 16574
rect 523052 16546 523908 16574
rect 527192 16546 527496 16574
rect 534092 16546 534580 16574
rect 484584 4820 484636 4826
rect 484584 4762 484636 4768
rect 481088 3528 481140 3534
rect 481088 3470 481140 3476
rect 481100 480 481128 3470
rect 484596 480 484624 4762
rect 488184 480 488212 16546
rect 491772 480 491800 16546
rect 495348 7608 495400 7614
rect 495348 7550 495400 7556
rect 495360 480 495388 7550
rect 498948 480 498976 16546
rect 502444 480 502472 16546
rect 506032 480 506060 16546
rect 509620 480 509648 16546
rect 513196 8968 513248 8974
rect 513196 8910 513248 8916
rect 513208 480 513236 8910
rect 516796 480 516824 16546
rect 520280 14476 520332 14482
rect 520280 14418 520332 14424
rect 520292 480 520320 14418
rect 523880 480 523908 16546
rect 527468 480 527496 16546
rect 531044 10328 531096 10334
rect 531044 10270 531096 10276
rect 531056 480 531084 10270
rect 534552 480 534580 16546
rect 536852 3534 536880 305594
rect 545120 304292 545172 304298
rect 545120 304234 545172 304240
rect 545132 16574 545160 304234
rect 547144 302932 547196 302938
rect 547144 302874 547196 302880
rect 545132 16546 545344 16574
rect 541716 15904 541768 15910
rect 541716 15846 541768 15852
rect 536840 3528 536892 3534
rect 536840 3470 536892 3476
rect 538128 3528 538180 3534
rect 538128 3470 538180 3476
rect 538140 480 538168 3470
rect 541728 480 541756 15846
rect 545316 480 545344 16546
rect 547156 4146 547184 302874
rect 554780 301504 554832 301510
rect 554780 301446 554832 301452
rect 552020 133204 552072 133210
rect 552020 133146 552072 133152
rect 552032 16574 552060 133146
rect 552032 16546 552428 16574
rect 547144 4140 547196 4146
rect 547144 4082 547196 4088
rect 548892 4140 548944 4146
rect 548892 4082 548944 4088
rect 548904 480 548932 4082
rect 552400 480 552428 16546
rect 554792 2922 554820 301446
rect 558196 3534 558224 318038
rect 563060 316736 563112 316742
rect 563060 316678 563112 316684
rect 563072 16574 563100 316678
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 565084 300144 565136 300150
rect 565084 300086 565136 300092
rect 563072 16546 563192 16574
rect 558184 3528 558236 3534
rect 558184 3470 558236 3476
rect 559564 3528 559616 3534
rect 559564 3470 559616 3476
rect 554780 2916 554832 2922
rect 554780 2858 554832 2864
rect 555976 2916 556028 2922
rect 555976 2858 556028 2864
rect 555988 480 556016 2858
rect 559576 480 559604 3470
rect 563164 480 563192 16546
rect 565096 3534 565124 300086
rect 567844 298784 567896 298790
rect 567844 298726 567896 298732
rect 567856 3534 567884 298726
rect 572720 297424 572772 297430
rect 572720 297366 572772 297372
rect 572732 16574 572760 297366
rect 576124 295996 576176 296002
rect 576124 295938 576176 295944
rect 572732 16546 573864 16574
rect 565084 3528 565136 3534
rect 565084 3470 565136 3476
rect 566740 3528 566792 3534
rect 566740 3470 566792 3476
rect 567844 3528 567896 3534
rect 567844 3470 567896 3476
rect 570236 3528 570288 3534
rect 570236 3470 570288 3476
rect 566752 480 566780 3470
rect 570248 480 570276 3470
rect 573836 480 573864 16546
rect 576136 4146 576164 295938
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 576124 4140 576176 4146
rect 576124 4082 576176 4088
rect 577412 4140 577464 4146
rect 577412 4082 577464 4088
rect 577424 480 577452 4082
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3514 653520 3570 653576
rect 3422 610408 3478 610464
rect 3330 553016 3386 553072
rect 3146 437960 3202 438016
rect 3146 423700 3202 423736
rect 3146 423680 3148 423700
rect 3148 423680 3200 423700
rect 3200 423680 3202 423700
rect 2962 366152 3018 366208
rect 3606 595992 3662 596048
rect 3790 538600 3846 538656
rect 3698 495488 3754 495544
rect 3606 380568 3662 380624
rect 3882 481072 3938 481128
rect 3238 323040 3294 323096
rect 3330 308760 3386 308816
rect 3146 280100 3148 280120
rect 3148 280100 3200 280120
rect 3200 280100 3202 280120
rect 3146 280064 3202 280100
rect 2870 265648 2926 265704
rect 3146 222536 3202 222592
rect 2870 193840 2926 193896
rect 3238 179424 3294 179480
rect 3146 150728 3202 150784
rect 3238 107616 3294 107672
rect 3330 64504 3386 64560
rect 3054 50088 3110 50144
rect 2870 21392 2926 21448
rect 3146 7112 3202 7168
rect 3514 236952 3570 237008
rect 3514 136312 3570 136368
rect 3514 93200 3570 93256
rect 321834 419056 321890 419112
rect 238022 418240 238078 418296
rect 237378 414704 237434 414760
rect 237378 408720 237434 408776
rect 237378 405748 237434 405784
rect 237378 405728 237380 405748
rect 237380 405728 237432 405748
rect 237432 405728 237434 405748
rect 237378 403028 237434 403064
rect 237378 403008 237380 403028
rect 237380 403008 237432 403028
rect 237432 403008 237434 403028
rect 237378 399200 237434 399256
rect 237378 396092 237434 396128
rect 237378 396072 237380 396092
rect 237380 396072 237432 396092
rect 237432 396072 237434 396092
rect 237378 390516 237434 390552
rect 237378 390496 237380 390516
rect 237380 390496 237432 390516
rect 237432 390496 237434 390516
rect 237378 387640 237434 387696
rect 237378 384956 237380 384976
rect 237380 384956 237432 384976
rect 237432 384956 237434 384976
rect 237378 384920 237434 384956
rect 237378 381792 237434 381848
rect 237378 377984 237434 378040
rect 237378 375300 237380 375320
rect 237380 375300 237432 375320
rect 237432 375300 237434 375320
rect 237378 375264 237434 375300
rect 237378 371456 237434 371512
rect 237378 365764 237434 365800
rect 237378 365744 237380 365764
rect 237380 365744 237432 365764
rect 237432 365744 237434 365764
rect 237378 358828 237434 358864
rect 237378 358808 237380 358828
rect 237380 358808 237432 358828
rect 237432 358808 237434 358828
rect 237378 352552 237434 352608
rect 237378 347692 237380 347712
rect 237380 347692 237432 347712
rect 237432 347692 237434 347712
rect 237378 347656 237434 347692
rect 237378 344528 237434 344584
rect 237378 340720 237434 340776
rect 237378 338036 237380 338056
rect 237380 338036 237432 338056
rect 237432 338036 237434 338056
rect 237378 338000 237434 338036
rect 237378 335144 237434 335200
rect 237378 332152 237434 332208
rect 321834 416336 321890 416392
rect 322202 413480 322258 413536
rect 238114 411576 238170 411632
rect 322202 410760 322258 410816
rect 322018 408040 322074 408096
rect 321834 405320 321890 405376
rect 322110 401648 322166 401704
rect 238298 393352 238354 393408
rect 238206 368464 238262 368520
rect 322754 398928 322810 398984
rect 322202 396480 322258 396536
rect 322478 394304 322534 394360
rect 321834 371728 321890 371784
rect 322478 391584 322534 391640
rect 322478 388864 322534 388920
rect 322478 386144 322534 386200
rect 322478 383424 322534 383480
rect 322478 380704 322534 380760
rect 322478 377984 322534 378040
rect 322294 374448 322350 374504
rect 321834 363432 321890 363488
rect 238298 361936 238354 361992
rect 321834 360712 321890 360768
rect 322662 368872 322718 368928
rect 322570 366152 322626 366208
rect 322478 357992 322534 358048
rect 238390 356088 238446 356144
rect 321650 355544 321706 355600
rect 322386 352552 322442 352608
rect 322018 349832 322074 349888
rect 238482 349424 238538 349480
rect 322018 347112 322074 347168
rect 322294 345092 322350 345128
rect 322294 345072 322296 345092
rect 322296 345072 322348 345092
rect 322348 345072 322350 345092
rect 322202 342216 322258 342272
rect 322294 339516 322350 339552
rect 322294 339496 322296 339516
rect 322296 339496 322348 339516
rect 322348 339496 322350 339516
rect 322202 336776 322258 336832
rect 322110 334056 322166 334112
rect 322110 331336 322166 331392
rect 580170 697992 580226 698048
rect 580262 686296 580318 686352
rect 580170 651072 580226 651128
rect 580170 604152 580226 604208
rect 579802 557232 579858 557288
rect 580170 545536 580226 545592
rect 579802 510312 579858 510368
rect 580170 498616 580226 498672
rect 579802 463392 579858 463448
rect 579618 416472 579674 416528
rect 580354 639376 580410 639432
rect 580446 592456 580502 592512
rect 580538 451696 580594 451752
rect 580630 404776 580686 404832
rect 580170 369552 580226 369608
rect 579986 357856 580042 357912
rect 580170 322632 580226 322688
rect 580170 310800 580226 310856
rect 580170 275712 580226 275768
rect 580170 263880 580226 263936
rect 579802 252184 579858 252240
rect 580170 228792 580226 228848
rect 580170 216960 580226 217016
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580257 686354 580323 686357
rect 583520 686354 584960 686444
rect 580257 686352 584960 686354
rect 580257 686296 580262 686352
rect 580318 686296 584960 686352
rect 580257 686294 584960 686296
rect 580257 686291 580323 686294
rect 583520 686204 584960 686294
rect -960 682124 480 682364
rect 583520 674508 584960 674748
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3509 653578 3575 653581
rect -960 653576 3575 653578
rect -960 653520 3514 653576
rect 3570 653520 3575 653576
rect -960 653518 3575 653520
rect -960 653428 480 653518
rect 3509 653515 3575 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580349 639434 580415 639437
rect 583520 639434 584960 639524
rect 580349 639432 584960 639434
rect 580349 639376 580354 639432
rect 580410 639376 584960 639432
rect 580349 639374 584960 639376
rect 580349 639371 580415 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 583520 627588 584960 627828
rect -960 624732 480 624972
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3601 596050 3667 596053
rect -960 596048 3667 596050
rect -960 595992 3606 596048
rect 3662 595992 3667 596048
rect -960 595990 3667 595992
rect -960 595900 480 595990
rect 3601 595987 3667 595990
rect 580441 592514 580507 592517
rect 583520 592514 584960 592604
rect 580441 592512 584960 592514
rect 580441 592456 580446 592512
rect 580502 592456 584960 592512
rect 580441 592454 584960 592456
rect 580441 592451 580507 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 583520 580668 584960 580908
rect 583520 568836 584960 569076
rect -960 567204 480 567444
rect 579797 557290 579863 557293
rect 583520 557290 584960 557380
rect 579797 557288 584960 557290
rect 579797 557232 579802 557288
rect 579858 557232 584960 557288
rect 579797 557230 584960 557232
rect 579797 557227 579863 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3325 553074 3391 553077
rect -960 553072 3391 553074
rect -960 553016 3330 553072
rect 3386 553016 3391 553072
rect -960 553014 3391 553016
rect -960 552924 480 553014
rect 3325 553011 3391 553014
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 3785 538658 3851 538661
rect -960 538656 3851 538658
rect -960 538600 3790 538656
rect 3846 538600 3851 538656
rect -960 538598 3851 538600
rect -960 538508 480 538598
rect 3785 538595 3851 538598
rect 583520 533748 584960 533988
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 579797 510370 579863 510373
rect 583520 510370 584960 510460
rect 579797 510368 584960 510370
rect 579797 510312 579802 510368
rect 579858 510312 584960 510368
rect 579797 510310 584960 510312
rect 579797 510307 579863 510310
rect 583520 510220 584960 510310
rect -960 509812 480 510052
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3693 495546 3759 495549
rect -960 495544 3759 495546
rect -960 495488 3698 495544
rect 3754 495488 3759 495544
rect -960 495486 3759 495488
rect -960 495396 480 495486
rect 3693 495483 3759 495486
rect 583520 486692 584960 486932
rect -960 481130 480 481220
rect 3877 481130 3943 481133
rect -960 481128 3943 481130
rect -960 481072 3882 481128
rect 3938 481072 3943 481128
rect -960 481070 3943 481072
rect -960 480980 480 481070
rect 3877 481067 3943 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 579797 463450 579863 463453
rect 583520 463450 584960 463540
rect 579797 463448 584960 463450
rect 579797 463392 579802 463448
rect 579858 463392 584960 463448
rect 579797 463390 584960 463392
rect 579797 463387 579863 463390
rect 583520 463300 584960 463390
rect -960 452284 480 452524
rect 580533 451754 580599 451757
rect 583520 451754 584960 451844
rect 580533 451752 584960 451754
rect 580533 451696 580538 451752
rect 580594 451696 584960 451752
rect 580533 451694 584960 451696
rect 580533 451691 580599 451694
rect 583520 451604 584960 451694
rect 583520 439772 584960 440012
rect -960 438018 480 438108
rect 3141 438018 3207 438021
rect -960 438016 3207 438018
rect -960 437960 3146 438016
rect 3202 437960 3207 438016
rect -960 437958 3207 437960
rect -960 437868 480 437958
rect 3141 437955 3207 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3141 423738 3207 423741
rect -960 423736 3207 423738
rect -960 423680 3146 423736
rect 3202 423680 3207 423736
rect -960 423678 3207 423680
rect -960 423588 480 423678
rect 3141 423675 3207 423678
rect 321829 419114 321895 419117
rect 319854 419112 321895 419114
rect 319854 419056 321834 419112
rect 321890 419056 321895 419112
rect 319854 419054 321895 419056
rect 319854 418608 319914 419054
rect 321829 419051 321895 419054
rect 238017 418298 238083 418301
rect 239998 418298 240058 418472
rect 238017 418296 240058 418298
rect 238017 418240 238022 418296
rect 238078 418240 240058 418296
rect 238017 418238 240058 418240
rect 238017 418235 238083 418238
rect 579613 416530 579679 416533
rect 583520 416530 584960 416620
rect 579613 416528 584960 416530
rect 579613 416472 579618 416528
rect 579674 416472 584960 416528
rect 579613 416470 584960 416472
rect 579613 416467 579679 416470
rect 321829 416394 321895 416397
rect 319854 416392 321895 416394
rect 319854 416336 321834 416392
rect 321890 416336 321895 416392
rect 583520 416380 584960 416470
rect 319854 416334 321895 416336
rect 319854 415888 319914 416334
rect 321829 416331 321895 416334
rect 237373 414762 237439 414765
rect 239998 414762 240058 415344
rect 237373 414760 240058 414762
rect 237373 414704 237378 414760
rect 237434 414704 240058 414760
rect 237373 414702 240058 414704
rect 237373 414699 237439 414702
rect 322197 413538 322263 413541
rect 319854 413536 322263 413538
rect 319854 413480 322202 413536
rect 322258 413480 322263 413536
rect 319854 413478 322263 413480
rect 319854 413168 319914 413478
rect 322197 413475 322263 413478
rect 238109 411634 238175 411637
rect 239998 411634 240058 412216
rect 238109 411632 240058 411634
rect 238109 411576 238114 411632
rect 238170 411576 240058 411632
rect 238109 411574 240058 411576
rect 238109 411571 238175 411574
rect 322197 410818 322263 410821
rect 319854 410816 322263 410818
rect 319854 410760 322202 410816
rect 322258 410760 322263 410816
rect 319854 410758 322263 410760
rect 319854 410448 319914 410758
rect 322197 410755 322263 410758
rect -960 409172 480 409412
rect 237373 408778 237439 408781
rect 239998 408778 240058 409088
rect 237373 408776 240058 408778
rect 237373 408720 237378 408776
rect 237434 408720 240058 408776
rect 237373 408718 240058 408720
rect 237373 408715 237439 408718
rect 322013 408098 322079 408101
rect 319854 408096 322079 408098
rect 319854 408040 322018 408096
rect 322074 408040 322079 408096
rect 319854 408038 322079 408040
rect 319854 407728 319914 408038
rect 322013 408035 322079 408038
rect 237373 405786 237439 405789
rect 239998 405786 240058 405960
rect 237373 405784 240058 405786
rect 237373 405728 237378 405784
rect 237434 405728 240058 405784
rect 237373 405726 240058 405728
rect 237373 405723 237439 405726
rect 321829 405378 321895 405381
rect 319854 405376 321895 405378
rect 319854 405320 321834 405376
rect 321890 405320 321895 405376
rect 319854 405318 321895 405320
rect 319854 405008 319914 405318
rect 321829 405315 321895 405318
rect 580625 404834 580691 404837
rect 583520 404834 584960 404924
rect 580625 404832 584960 404834
rect 580625 404776 580630 404832
rect 580686 404776 584960 404832
rect 580625 404774 584960 404776
rect 580625 404771 580691 404774
rect 583520 404684 584960 404774
rect 237373 403066 237439 403069
rect 237373 403064 240058 403066
rect 237373 403008 237378 403064
rect 237434 403008 240058 403064
rect 237373 403006 240058 403008
rect 237373 403003 237439 403006
rect 239998 402968 240058 403006
rect 319854 401706 319914 402288
rect 322105 401706 322171 401709
rect 319854 401704 322171 401706
rect 319854 401648 322110 401704
rect 322166 401648 322171 401704
rect 319854 401646 322171 401648
rect 322105 401643 322171 401646
rect 237373 399258 237439 399261
rect 239998 399258 240058 399840
rect 237373 399256 240058 399258
rect 237373 399200 237378 399256
rect 237434 399200 240058 399256
rect 237373 399198 240058 399200
rect 237373 399195 237439 399198
rect 319854 398986 319914 399568
rect 322749 398986 322815 398989
rect 319854 398984 322815 398986
rect 319854 398928 322754 398984
rect 322810 398928 322815 398984
rect 319854 398926 322815 398928
rect 322749 398923 322815 398926
rect 237373 396130 237439 396133
rect 239998 396130 240058 396712
rect 319854 396538 319914 396848
rect 322197 396538 322263 396541
rect 319854 396536 322263 396538
rect 319854 396480 322202 396536
rect 322258 396480 322263 396536
rect 319854 396478 322263 396480
rect 322197 396475 322263 396478
rect 237373 396128 240058 396130
rect 237373 396072 237378 396128
rect 237434 396072 240058 396128
rect 237373 396070 240058 396072
rect 237373 396067 237439 396070
rect -960 394892 480 395132
rect 322473 394362 322539 394365
rect 319854 394360 322539 394362
rect 319854 394304 322478 394360
rect 322534 394304 322539 394360
rect 319854 394302 322539 394304
rect 319854 394128 319914 394302
rect 322473 394299 322539 394302
rect 238293 393410 238359 393413
rect 239998 393410 240058 393584
rect 238293 393408 240058 393410
rect 238293 393352 238298 393408
rect 238354 393352 240058 393408
rect 238293 393350 240058 393352
rect 238293 393347 238359 393350
rect 583520 392852 584960 393092
rect 322473 391642 322539 391645
rect 319854 391640 322539 391642
rect 319854 391584 322478 391640
rect 322534 391584 322539 391640
rect 319854 391582 322539 391584
rect 319854 391408 319914 391582
rect 322473 391579 322539 391582
rect 237373 390554 237439 390557
rect 237373 390552 240058 390554
rect 237373 390496 237378 390552
rect 237434 390496 240058 390552
rect 237373 390494 240058 390496
rect 237373 390491 237439 390494
rect 239998 390456 240058 390494
rect 322473 388922 322539 388925
rect 319854 388920 322539 388922
rect 319854 388864 322478 388920
rect 322534 388864 322539 388920
rect 319854 388862 322539 388864
rect 319854 388688 319914 388862
rect 322473 388859 322539 388862
rect 237373 387698 237439 387701
rect 237373 387696 240058 387698
rect 237373 387640 237378 387696
rect 237434 387640 240058 387696
rect 237373 387638 240058 387640
rect 237373 387635 237439 387638
rect 239998 387328 240058 387638
rect 322473 386202 322539 386205
rect 319854 386200 322539 386202
rect 319854 386144 322478 386200
rect 322534 386144 322539 386200
rect 319854 386142 322539 386144
rect 319854 385968 319914 386142
rect 322473 386139 322539 386142
rect 237373 384978 237439 384981
rect 237373 384976 240058 384978
rect 237373 384920 237378 384976
rect 237434 384920 240058 384976
rect 237373 384918 240058 384920
rect 237373 384915 237439 384918
rect 239998 384336 240058 384918
rect 322473 383482 322539 383485
rect 319854 383480 322539 383482
rect 319854 383424 322478 383480
rect 322534 383424 322539 383480
rect 319854 383422 322539 383424
rect 319854 383248 319914 383422
rect 322473 383419 322539 383422
rect 237373 381850 237439 381853
rect 237373 381848 240058 381850
rect 237373 381792 237378 381848
rect 237434 381792 240058 381848
rect 237373 381790 240058 381792
rect 237373 381787 237439 381790
rect 239998 381208 240058 381790
rect 583520 381156 584960 381396
rect 322473 380762 322539 380765
rect 319854 380760 322539 380762
rect -960 380626 480 380716
rect 319854 380704 322478 380760
rect 322534 380704 322539 380760
rect 319854 380702 322539 380704
rect 3601 380626 3667 380629
rect -960 380624 3667 380626
rect -960 380568 3606 380624
rect 3662 380568 3667 380624
rect -960 380566 3667 380568
rect -960 380476 480 380566
rect 3601 380563 3667 380566
rect 319854 380528 319914 380702
rect 322473 380699 322539 380702
rect 237373 378042 237439 378045
rect 239998 378042 240058 378080
rect 322473 378042 322539 378045
rect 237373 378040 240058 378042
rect 237373 377984 237378 378040
rect 237434 377984 240058 378040
rect 237373 377982 240058 377984
rect 319854 378040 322539 378042
rect 319854 377984 322478 378040
rect 322534 377984 322539 378040
rect 319854 377982 322539 377984
rect 237373 377979 237439 377982
rect 319854 377808 319914 377982
rect 322473 377979 322539 377982
rect 237373 375322 237439 375325
rect 237373 375320 240058 375322
rect 237373 375264 237378 375320
rect 237434 375264 240058 375320
rect 237373 375262 240058 375264
rect 237373 375259 237439 375262
rect 239998 374952 240058 375262
rect 319854 374506 319914 374952
rect 322289 374506 322355 374509
rect 319854 374504 322355 374506
rect 319854 374448 322294 374504
rect 322350 374448 322355 374504
rect 319854 374446 322355 374448
rect 322289 374443 322355 374446
rect 237373 371514 237439 371517
rect 239998 371514 240058 371824
rect 319854 371786 319914 372232
rect 321829 371786 321895 371789
rect 319854 371784 321895 371786
rect 319854 371728 321834 371784
rect 321890 371728 321895 371784
rect 319854 371726 321895 371728
rect 321829 371723 321895 371726
rect 237373 371512 240058 371514
rect 237373 371456 237378 371512
rect 237434 371456 240058 371512
rect 237373 371454 240058 371456
rect 237373 371451 237439 371454
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 319854 368930 319914 369512
rect 583520 369460 584960 369550
rect 322657 368930 322723 368933
rect 319854 368928 322723 368930
rect 319854 368872 322662 368928
rect 322718 368872 322723 368928
rect 319854 368870 322723 368872
rect 322657 368867 322723 368870
rect 238201 368522 238267 368525
rect 239998 368522 240058 368696
rect 238201 368520 240058 368522
rect 238201 368464 238206 368520
rect 238262 368464 240058 368520
rect 238201 368462 240058 368464
rect 238201 368459 238267 368462
rect -960 366210 480 366300
rect 2957 366210 3023 366213
rect -960 366208 3023 366210
rect -960 366152 2962 366208
rect 3018 366152 3023 366208
rect -960 366150 3023 366152
rect 319854 366210 319914 366792
rect 322565 366210 322631 366213
rect 319854 366208 322631 366210
rect 319854 366152 322570 366208
rect 322626 366152 322631 366208
rect 319854 366150 322631 366152
rect -960 366060 480 366150
rect 2957 366147 3023 366150
rect 322565 366147 322631 366150
rect 237373 365802 237439 365805
rect 237373 365800 240058 365802
rect 237373 365744 237378 365800
rect 237434 365744 240058 365800
rect 237373 365742 240058 365744
rect 237373 365739 237439 365742
rect 239998 365704 240058 365742
rect 319854 363490 319914 364072
rect 321829 363490 321895 363493
rect 319854 363488 321895 363490
rect 319854 363432 321834 363488
rect 321890 363432 321895 363488
rect 319854 363430 321895 363432
rect 321829 363427 321895 363430
rect 238293 361994 238359 361997
rect 239998 361994 240058 362576
rect 238293 361992 240058 361994
rect 238293 361936 238298 361992
rect 238354 361936 240058 361992
rect 238293 361934 240058 361936
rect 238293 361931 238359 361934
rect 319854 360770 319914 361352
rect 321829 360770 321895 360773
rect 319854 360768 321895 360770
rect 319854 360712 321834 360768
rect 321890 360712 321895 360768
rect 319854 360710 321895 360712
rect 321829 360707 321895 360710
rect 237373 358866 237439 358869
rect 239998 358866 240058 359448
rect 237373 358864 240058 358866
rect 237373 358808 237378 358864
rect 237434 358808 240058 358864
rect 237373 358806 240058 358808
rect 237373 358803 237439 358806
rect 319854 358050 319914 358632
rect 322473 358050 322539 358053
rect 319854 358048 322539 358050
rect 319854 357992 322478 358048
rect 322534 357992 322539 358048
rect 319854 357990 322539 357992
rect 322473 357987 322539 357990
rect 579981 357914 580047 357917
rect 583520 357914 584960 358004
rect 579981 357912 584960 357914
rect 579981 357856 579986 357912
rect 580042 357856 584960 357912
rect 579981 357854 584960 357856
rect 579981 357851 580047 357854
rect 583520 357764 584960 357854
rect 238385 356146 238451 356149
rect 239998 356146 240058 356320
rect 238385 356144 240058 356146
rect 238385 356088 238390 356144
rect 238446 356088 240058 356144
rect 238385 356086 240058 356088
rect 238385 356083 238451 356086
rect 319854 355602 319914 355912
rect 321645 355602 321711 355605
rect 319854 355600 321711 355602
rect 319854 355544 321650 355600
rect 321706 355544 321711 355600
rect 319854 355542 321711 355544
rect 321645 355539 321711 355542
rect 237373 352610 237439 352613
rect 239998 352610 240058 353192
rect 237373 352608 240058 352610
rect 237373 352552 237378 352608
rect 237434 352552 240058 352608
rect 237373 352550 240058 352552
rect 319854 352610 319914 353192
rect 322381 352610 322447 352613
rect 319854 352608 322447 352610
rect 319854 352552 322386 352608
rect 322442 352552 322447 352608
rect 319854 352550 322447 352552
rect 237373 352547 237439 352550
rect 322381 352547 322447 352550
rect -960 351780 480 352020
rect 238477 349482 238543 349485
rect 239998 349482 240058 350064
rect 319854 349890 319914 350472
rect 322013 349890 322079 349893
rect 319854 349888 322079 349890
rect 319854 349832 322018 349888
rect 322074 349832 322079 349888
rect 319854 349830 322079 349832
rect 322013 349827 322079 349830
rect 238477 349480 240058 349482
rect 238477 349424 238482 349480
rect 238538 349424 240058 349480
rect 238477 349422 240058 349424
rect 238477 349419 238543 349422
rect 237373 347714 237439 347717
rect 237373 347712 240058 347714
rect 237373 347656 237378 347712
rect 237434 347656 240058 347712
rect 237373 347654 240058 347656
rect 237373 347651 237439 347654
rect 239998 347072 240058 347654
rect 319854 347170 319914 347752
rect 322013 347170 322079 347173
rect 319854 347168 322079 347170
rect 319854 347112 322018 347168
rect 322074 347112 322079 347168
rect 319854 347110 322079 347112
rect 322013 347107 322079 347110
rect 583520 345932 584960 346172
rect 322289 345130 322355 345133
rect 319854 345128 322355 345130
rect 319854 345072 322294 345128
rect 322350 345072 322355 345128
rect 319854 345070 322355 345072
rect 319854 345032 319914 345070
rect 322289 345067 322355 345070
rect 237373 344586 237439 344589
rect 237373 344584 240058 344586
rect 237373 344528 237378 344584
rect 237434 344528 240058 344584
rect 237373 344526 240058 344528
rect 237373 344523 237439 344526
rect 239998 343944 240058 344526
rect 319854 342274 319914 342312
rect 322197 342274 322263 342277
rect 319854 342272 322263 342274
rect 319854 342216 322202 342272
rect 322258 342216 322263 342272
rect 319854 342214 322263 342216
rect 322197 342211 322263 342214
rect 237373 340778 237439 340781
rect 239998 340778 240058 340816
rect 237373 340776 240058 340778
rect 237373 340720 237378 340776
rect 237434 340720 240058 340776
rect 237373 340718 240058 340720
rect 237373 340715 237439 340718
rect 319854 339554 319914 339592
rect 322289 339554 322355 339557
rect 319854 339552 322355 339554
rect 319854 339496 322294 339552
rect 322350 339496 322355 339552
rect 319854 339494 322355 339496
rect 322289 339491 322355 339494
rect 237373 338058 237439 338061
rect 237373 338056 240058 338058
rect 237373 338000 237378 338056
rect 237434 338000 240058 338056
rect 237373 337998 240058 338000
rect 237373 337995 237439 337998
rect 239998 337688 240058 337998
rect -960 337364 480 337604
rect 319854 336834 319914 336872
rect 322197 336834 322263 336837
rect 319854 336832 322263 336834
rect 319854 336776 322202 336832
rect 322258 336776 322263 336832
rect 319854 336774 322263 336776
rect 322197 336771 322263 336774
rect 237373 335202 237439 335205
rect 237373 335200 240058 335202
rect 237373 335144 237378 335200
rect 237434 335144 240058 335200
rect 237373 335142 240058 335144
rect 237373 335139 237439 335142
rect 239998 334560 240058 335142
rect 583520 334236 584960 334476
rect 319854 334114 319914 334152
rect 322105 334114 322171 334117
rect 319854 334112 322171 334114
rect 319854 334056 322110 334112
rect 322166 334056 322171 334112
rect 319854 334054 322171 334056
rect 322105 334051 322171 334054
rect 237373 332210 237439 332213
rect 237373 332208 240058 332210
rect 237373 332152 237378 332208
rect 237434 332152 240058 332208
rect 237373 332150 240058 332152
rect 237373 332147 237439 332150
rect 239998 331568 240058 332150
rect 319854 331394 319914 331432
rect 322105 331394 322171 331397
rect 319854 331392 322171 331394
rect 319854 331336 322110 331392
rect 322166 331336 322171 331392
rect 319854 331334 322171 331336
rect 322105 331331 322171 331334
rect -960 323098 480 323188
rect 3233 323098 3299 323101
rect -960 323096 3299 323098
rect -960 323040 3238 323096
rect 3294 323040 3299 323096
rect -960 323038 3299 323040
rect -960 322948 480 323038
rect 3233 323035 3299 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 583520 299012 584960 299252
rect -960 294252 480 294492
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3141 280122 3207 280125
rect -960 280120 3207 280122
rect -960 280064 3146 280120
rect 3202 280064 3207 280120
rect -960 280062 3207 280064
rect -960 279972 480 280062
rect 3141 280059 3207 280062
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect -960 265706 480 265796
rect 2865 265706 2931 265709
rect -960 265704 2931 265706
rect -960 265648 2870 265704
rect 2926 265648 2931 265704
rect -960 265646 2931 265648
rect -960 265556 480 265646
rect 2865 265643 2931 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251140 480 251380
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3509 237010 3575 237013
rect -960 237008 3575 237010
rect -960 236952 3514 237008
rect 3570 236952 3575 237008
rect -960 236950 3575 236952
rect -960 236860 480 236950
rect 3509 236947 3575 236950
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect -960 208028 480 208268
rect 583520 205172 584960 205412
rect -960 193898 480 193988
rect 2865 193898 2931 193901
rect -960 193896 2931 193898
rect -960 193840 2870 193896
rect 2926 193840 2931 193896
rect -960 193838 2931 193840
rect -960 193748 480 193838
rect 2865 193835 2931 193838
rect 583520 193476 584960 193716
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect -960 164916 480 165156
rect 583520 158252 584960 158492
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 583520 146556 584960 146796
rect -960 136370 480 136460
rect 3509 136370 3575 136373
rect -960 136368 3575 136370
rect -960 136312 3514 136368
rect 3570 136312 3575 136368
rect -960 136310 3575 136312
rect -960 136220 480 136310
rect 3509 136307 3575 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 121940 480 122180
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 583520 99636 584960 99876
rect -960 93258 480 93348
rect 3509 93258 3575 93261
rect -960 93256 3575 93258
rect -960 93200 3514 93256
rect 3570 93200 3575 93256
rect -960 93198 3575 93200
rect -960 93108 480 93198
rect 3509 93195 3575 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect -960 78828 480 79068
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3049 50146 3115 50149
rect -960 50144 3115 50146
rect -960 50088 3054 50144
rect 3110 50088 3115 50144
rect -960 50086 3115 50088
rect -960 49996 480 50086
rect 3049 50083 3115 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35716 480 35956
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect -960 21450 480 21540
rect 2865 21450 2931 21453
rect -960 21448 2931 21450
rect -960 21392 2870 21448
rect 2926 21392 2931 21448
rect -960 21390 2931 21392
rect -960 21300 480 21390
rect 2865 21387 2931 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3141 7170 3207 7173
rect -960 7168 3207 7170
rect -960 7112 3146 7168
rect 3202 7112 3207 7168
rect -960 7110 3207 7112
rect -960 7020 480 7110
rect 3141 7107 3207 7110
rect 583520 5796 584960 6036
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 421000 239004 455498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 421000 242604 423098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 421000 246204 426698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 421000 253404 433898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 421000 257004 437498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 421000 260604 441098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 421000 264204 444698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 421000 271404 451898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 421000 275004 455498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 421000 278604 423098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 421000 282204 426698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 421000 289404 433898
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 421000 293004 437498
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 421000 296604 441098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 421000 300204 444698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 421000 307404 451898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 421000 311004 455498
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 421000 314604 423098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 421000 318204 426698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 259568 416454 259888 416476
rect 259568 416218 259610 416454
rect 259846 416218 259888 416454
rect 259568 416134 259888 416218
rect 259568 415898 259610 416134
rect 259846 415898 259888 416134
rect 259568 415876 259888 415898
rect 290288 416454 290608 416476
rect 290288 416218 290330 416454
rect 290566 416218 290608 416454
rect 290288 416134 290608 416218
rect 290288 415898 290330 416134
rect 290566 415898 290608 416134
rect 290288 415876 290608 415898
rect 244208 398454 244528 398476
rect 244208 398218 244250 398454
rect 244486 398218 244528 398454
rect 244208 398134 244528 398218
rect 244208 397898 244250 398134
rect 244486 397898 244528 398134
rect 244208 397876 244528 397898
rect 274928 398454 275248 398476
rect 274928 398218 274970 398454
rect 275206 398218 275248 398454
rect 274928 398134 275248 398218
rect 274928 397898 274970 398134
rect 275206 397898 275248 398134
rect 274928 397876 275248 397898
rect 305648 398454 305968 398476
rect 305648 398218 305690 398454
rect 305926 398218 305968 398454
rect 305648 398134 305968 398218
rect 305648 397898 305690 398134
rect 305926 397898 305968 398134
rect 305648 397876 305968 397898
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 259568 380454 259888 380476
rect 259568 380218 259610 380454
rect 259846 380218 259888 380454
rect 259568 380134 259888 380218
rect 259568 379898 259610 380134
rect 259846 379898 259888 380134
rect 259568 379876 259888 379898
rect 290288 380454 290608 380476
rect 290288 380218 290330 380454
rect 290566 380218 290608 380454
rect 290288 380134 290608 380218
rect 290288 379898 290330 380134
rect 290566 379898 290608 380134
rect 290288 379876 290608 379898
rect 244208 362454 244528 362476
rect 244208 362218 244250 362454
rect 244486 362218 244528 362454
rect 244208 362134 244528 362218
rect 244208 361898 244250 362134
rect 244486 361898 244528 362134
rect 244208 361876 244528 361898
rect 274928 362454 275248 362476
rect 274928 362218 274970 362454
rect 275206 362218 275248 362454
rect 274928 362134 275248 362218
rect 274928 361898 274970 362134
rect 275206 361898 275248 362134
rect 274928 361876 275248 361898
rect 305648 362454 305968 362476
rect 305648 362218 305690 362454
rect 305926 362218 305968 362454
rect 305648 362134 305968 362218
rect 305648 361898 305690 362134
rect 305926 361898 305968 362134
rect 305648 361876 305968 361898
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 259568 344454 259888 344476
rect 259568 344218 259610 344454
rect 259846 344218 259888 344454
rect 259568 344134 259888 344218
rect 259568 343898 259610 344134
rect 259846 343898 259888 344134
rect 259568 343876 259888 343898
rect 290288 344454 290608 344476
rect 290288 344218 290330 344454
rect 290566 344218 290608 344454
rect 290288 344134 290608 344218
rect 290288 343898 290330 344134
rect 290566 343898 290608 344134
rect 290288 343876 290608 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 312054 239004 329000
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 315654 242604 329000
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 319254 246204 329000
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 326454 253404 329000
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 294054 257004 329000
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 297654 260604 329000
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 301254 264204 329000
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 308454 271404 329000
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 312054 275004 329000
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 315654 278604 329000
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 319254 282204 329000
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 326454 289404 329000
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 294054 293004 329000
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 297654 296604 329000
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 301254 300204 329000
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 308454 307404 329000
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 312054 311004 329000
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 315654 314604 329000
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 319254 318204 329000
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 259610 416218 259846 416454
rect 259610 415898 259846 416134
rect 290330 416218 290566 416454
rect 290330 415898 290566 416134
rect 244250 398218 244486 398454
rect 244250 397898 244486 398134
rect 274970 398218 275206 398454
rect 274970 397898 275206 398134
rect 305690 398218 305926 398454
rect 305690 397898 305926 398134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 259610 380218 259846 380454
rect 259610 379898 259846 380134
rect 290330 380218 290566 380454
rect 290330 379898 290566 380134
rect 244250 362218 244486 362454
rect 244250 361898 244486 362134
rect 274970 362218 275206 362454
rect 274970 361898 275206 362134
rect 305690 362218 305926 362454
rect 305690 361898 305926 362134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 259610 344218 259846 344454
rect 259610 343898 259846 344134
rect 290330 344218 290566 344454
rect 290330 343898 290566 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 259568 416476 259888 416478
rect 290288 416476 290608 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 259610 416454
rect 259846 416218 290330 416454
rect 290566 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 259610 416134
rect 259846 415898 290330 416134
rect 290566 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 259568 415874 259888 415876
rect 290288 415874 290608 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 244208 398476 244528 398478
rect 274928 398476 275248 398478
rect 305648 398476 305968 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 244250 398454
rect 244486 398218 274970 398454
rect 275206 398218 305690 398454
rect 305926 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 244250 398134
rect 244486 397898 274970 398134
rect 275206 397898 305690 398134
rect 305926 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 244208 397874 244528 397876
rect 274928 397874 275248 397876
rect 305648 397874 305968 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 259568 380476 259888 380478
rect 290288 380476 290608 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 259610 380454
rect 259846 380218 290330 380454
rect 290566 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 259610 380134
rect 259846 379898 290330 380134
rect 290566 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 259568 379874 259888 379876
rect 290288 379874 290608 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 244208 362476 244528 362478
rect 274928 362476 275248 362478
rect 305648 362476 305968 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 244250 362454
rect 244486 362218 274970 362454
rect 275206 362218 305690 362454
rect 305926 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 244250 362134
rect 244486 361898 274970 362134
rect 275206 361898 305690 362134
rect 305926 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 244208 361874 244528 361876
rect 274928 361874 275248 361876
rect 305648 361874 305968 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 259568 344476 259888 344478
rect 290288 344476 290608 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 259610 344454
rect 259846 344218 290330 344454
rect 290566 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 259610 344134
rect 259846 343898 290330 344134
rect 290566 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 259568 343874 259888 343876
rect 290288 343874 290608 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use user_proj_top  user_proj_top
timestamp 1612364373
transform 1 0 240000 0 1 330000
box 0 0 80000 90000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew signal input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew signal input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew signal input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew signal input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew signal input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew signal input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew signal input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew signal input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew signal input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew signal input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew signal input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew signal input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew signal input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew signal input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew signal input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew signal input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew signal input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew signal input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew signal input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew signal input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew signal input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew signal input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew signal input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew signal input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew signal input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew signal input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew signal input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew signal input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew signal input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew signal tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew signal tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew signal tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew signal tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew signal tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew signal tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew signal tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew signal tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew signal tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew signal tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew signal tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew signal tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew signal tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew signal tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew signal tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew signal tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew signal tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew signal tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew signal tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew signal tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew signal tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew signal tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew signal tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew signal tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew signal tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew signal tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew signal tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew signal tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew signal tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew signal tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew signal tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew signal tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew signal tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew signal tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew signal tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew signal tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew signal tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew signal tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew signal tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew signal tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew signal tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew signal tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew signal tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew signal tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew signal tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew signal tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew signal tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew signal tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew signal tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew signal tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew signal tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew signal tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew signal tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew signal tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew signal tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew signal tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew signal tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew signal tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew signal tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew signal tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew signal tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew signal tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew signal tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew signal tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew signal tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew signal tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew signal tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew signal tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew signal tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew signal tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew signal tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew signal tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew signal tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew signal tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew signal tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew signal tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew signal tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew signal tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew signal tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew signal tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew signal tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew signal tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew signal tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew signal tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew signal tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew signal tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew signal tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew signal tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew signal tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew signal tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew signal tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew signal tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew signal tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew signal tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew signal tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew signal tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew signal tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew signal tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew signal tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew signal tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew signal tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew signal tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew signal tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew signal tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew signal tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew signal tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew signal tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew signal tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew signal tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew signal tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew signal tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew signal tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew signal tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew signal tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew signal tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew signal tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew signal tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew signal tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew signal tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew signal tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew signal tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew signal tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew signal tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew signal tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew signal tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew signal tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew signal tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew signal tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew signal tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew signal tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew signal tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew signal tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew signal tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew signal tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew signal tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew signal tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew signal tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew signal tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew signal tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew signal tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew signal tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew signal tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew signal tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew signal tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew signal tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew signal tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew signal tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew signal tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew signal tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew signal tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew signal tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew signal tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew signal tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew signal tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew signal tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew signal tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew signal tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew signal tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew signal tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew signal tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew signal tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew signal tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew signal tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew signal tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew signal tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew signal tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew signal tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew signal tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew signal tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew signal tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew signal tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew signal tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew signal tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew signal tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew signal tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew signal tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew signal tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew signal tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew signal tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew signal tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew signal tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew signal tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew signal tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew signal tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew signal tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew signal input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew signal input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew signal input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew signal input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew signal input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew signal input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew signal input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew signal input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew signal input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew signal input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew signal input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew signal input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew signal input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew signal input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew signal input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew signal input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew signal input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew signal input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew signal input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew signal input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew signal input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew signal input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew signal input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew signal input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew signal input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew signal input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew signal input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew signal input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew signal input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew signal input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew signal input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew signal input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew signal input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew signal input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew signal input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew signal input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew signal input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew signal input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew signal input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew signal input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew signal input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew signal input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew signal input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew signal input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew signal input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew signal input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew signal input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew signal input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew signal input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew signal input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew signal input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew signal input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew signal input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew signal input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew signal input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew signal input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew signal input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew signal input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew signal input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew signal input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew signal input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew signal input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew signal input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew signal input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew signal input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew signal input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew signal input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew signal input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew signal input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew signal input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew signal input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew signal input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew signal input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew signal input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew signal input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew signal input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew signal input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew signal input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew signal input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew signal input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew signal input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew signal input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew signal input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew signal input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew signal input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew signal input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew signal input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew signal input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew signal input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew signal input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew signal input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew signal input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew signal input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew signal input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew signal input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew signal input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew signal input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew signal input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew signal input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew signal input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew signal input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew signal input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew signal input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew signal input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew signal input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew signal input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew signal input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew signal input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew signal input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew signal input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew signal input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew signal input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew signal input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew signal input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew signal input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew signal input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew signal input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew signal input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew signal input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew signal input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew signal input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew signal input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew signal input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew signal input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew signal input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew signal input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew signal input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew signal input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew signal input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew signal input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew signal input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew signal input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew signal input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew signal input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew signal input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew signal input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew signal input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew signal input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew signal input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew signal input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew signal input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew signal input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew signal input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew signal input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew signal input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew signal input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew signal input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew signal input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew signal input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew signal input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew signal input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew signal input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew signal input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew signal input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew signal input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew signal input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew signal input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew signal input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew signal input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew signal input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew signal input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew signal input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew signal input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew signal input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew signal input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew signal input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew signal input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew signal input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew signal input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew signal input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew signal input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew signal input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew signal input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew signal input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew signal input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew signal input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew signal input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew signal input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew signal input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew signal input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew signal input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew signal input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew signal input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew signal input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew signal input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew signal input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew signal input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew signal input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew signal tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew signal tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew signal tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew signal tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew signal tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew signal tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew signal tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew signal tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew signal tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew signal tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew signal tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew signal tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew signal tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew signal tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew signal tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew signal tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew signal tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew signal tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew signal tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew signal tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew signal tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew signal tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew signal tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew signal tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew signal tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew signal tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew signal tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew signal tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew signal tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew signal tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew signal tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew signal tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew signal input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew signal input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew signal input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew signal input
rlabel metal4 s 576804 -1864 577404 705800 6 vccd1
port 636 nsew power bidirectional
rlabel metal4 s 540804 -1864 541404 705800 6 vccd1
port 637 nsew power bidirectional
rlabel metal4 s 504804 -1864 505404 705800 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 468804 -1864 469404 705800 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 432804 -1864 433404 705800 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 396804 -1864 397404 705800 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 360804 -1864 361404 705800 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 324804 -1864 325404 705800 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 288804 421000 289404 705800 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 252804 421000 253404 705800 6 vccd1
port 645 nsew power bidirectional
rlabel metal4 s 216804 -1864 217404 705800 6 vccd1
port 646 nsew power bidirectional
rlabel metal4 s 180804 -1864 181404 705800 6 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 144804 -1864 145404 705800 6 vccd1
port 648 nsew power bidirectional
rlabel metal4 s 108804 -1864 109404 705800 6 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 72804 -1864 73404 705800 6 vccd1
port 650 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 705800 6 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 705800 6 vccd1
port 652 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 653 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 654 nsew power bidirectional
rlabel metal4 s 288804 -1864 289404 329000 6 vccd1
port 655 nsew power bidirectional
rlabel metal4 s 252804 -1864 253404 329000 6 vccd1
port 656 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1
port 657 nsew power bidirectional
rlabel metal5 s -2936 685876 586860 686476 6 vccd1
port 658 nsew power bidirectional
rlabel metal5 s -2936 649876 586860 650476 6 vccd1
port 659 nsew power bidirectional
rlabel metal5 s -2936 613876 586860 614476 6 vccd1
port 660 nsew power bidirectional
rlabel metal5 s -2936 577876 586860 578476 6 vccd1
port 661 nsew power bidirectional
rlabel metal5 s -2936 541876 586860 542476 6 vccd1
port 662 nsew power bidirectional
rlabel metal5 s -2936 505876 586860 506476 6 vccd1
port 663 nsew power bidirectional
rlabel metal5 s -2936 469876 586860 470476 6 vccd1
port 664 nsew power bidirectional
rlabel metal5 s -2936 433876 586860 434476 6 vccd1
port 665 nsew power bidirectional
rlabel metal5 s -2936 397876 586860 398476 6 vccd1
port 666 nsew power bidirectional
rlabel metal5 s -2936 361876 586860 362476 6 vccd1
port 667 nsew power bidirectional
rlabel metal5 s -2936 325876 586860 326476 6 vccd1
port 668 nsew power bidirectional
rlabel metal5 s -2936 289876 586860 290476 6 vccd1
port 669 nsew power bidirectional
rlabel metal5 s -2936 253876 586860 254476 6 vccd1
port 670 nsew power bidirectional
rlabel metal5 s -2936 217876 586860 218476 6 vccd1
port 671 nsew power bidirectional
rlabel metal5 s -2936 181876 586860 182476 6 vccd1
port 672 nsew power bidirectional
rlabel metal5 s -2936 145876 586860 146476 6 vccd1
port 673 nsew power bidirectional
rlabel metal5 s -2936 109876 586860 110476 6 vccd1
port 674 nsew power bidirectional
rlabel metal5 s -2936 73876 586860 74476 6 vccd1
port 675 nsew power bidirectional
rlabel metal5 s -2936 37876 586860 38476 6 vccd1
port 676 nsew power bidirectional
rlabel metal5 s -2936 1876 586860 2476 6 vccd1
port 677 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 678 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 679 nsew ground bidirectional
rlabel metal4 s 558804 -1864 559404 705800 6 vssd1
port 680 nsew ground bidirectional
rlabel metal4 s 522804 -1864 523404 705800 6 vssd1
port 681 nsew ground bidirectional
rlabel metal4 s 486804 -1864 487404 705800 6 vssd1
port 682 nsew ground bidirectional
rlabel metal4 s 450804 -1864 451404 705800 6 vssd1
port 683 nsew ground bidirectional
rlabel metal4 s 414804 -1864 415404 705800 6 vssd1
port 684 nsew ground bidirectional
rlabel metal4 s 378804 -1864 379404 705800 6 vssd1
port 685 nsew ground bidirectional
rlabel metal4 s 342804 -1864 343404 705800 6 vssd1
port 686 nsew ground bidirectional
rlabel metal4 s 306804 421000 307404 705800 6 vssd1
port 687 nsew ground bidirectional
rlabel metal4 s 270804 421000 271404 705800 6 vssd1
port 688 nsew ground bidirectional
rlabel metal4 s 234804 -1864 235404 705800 6 vssd1
port 689 nsew ground bidirectional
rlabel metal4 s 198804 -1864 199404 705800 6 vssd1
port 690 nsew ground bidirectional
rlabel metal4 s 162804 -1864 163404 705800 6 vssd1
port 691 nsew ground bidirectional
rlabel metal4 s 126804 -1864 127404 705800 6 vssd1
port 692 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 705800 6 vssd1
port 693 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 705800 6 vssd1
port 694 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 705800 6 vssd1
port 695 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 696 nsew ground bidirectional
rlabel metal4 s 306804 -1864 307404 329000 6 vssd1
port 697 nsew ground bidirectional
rlabel metal4 s 270804 -1864 271404 329000 6 vssd1
port 698 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1
port 699 nsew ground bidirectional
rlabel metal5 s -2936 667876 586860 668476 6 vssd1
port 700 nsew ground bidirectional
rlabel metal5 s -2936 631876 586860 632476 6 vssd1
port 701 nsew ground bidirectional
rlabel metal5 s -2936 595876 586860 596476 6 vssd1
port 702 nsew ground bidirectional
rlabel metal5 s -2936 559876 586860 560476 6 vssd1
port 703 nsew ground bidirectional
rlabel metal5 s -2936 523876 586860 524476 6 vssd1
port 704 nsew ground bidirectional
rlabel metal5 s -2936 487876 586860 488476 6 vssd1
port 705 nsew ground bidirectional
rlabel metal5 s -2936 451876 586860 452476 6 vssd1
port 706 nsew ground bidirectional
rlabel metal5 s -2936 415876 586860 416476 6 vssd1
port 707 nsew ground bidirectional
rlabel metal5 s -2936 379876 586860 380476 6 vssd1
port 708 nsew ground bidirectional
rlabel metal5 s -2936 343876 586860 344476 6 vssd1
port 709 nsew ground bidirectional
rlabel metal5 s -2936 307876 586860 308476 6 vssd1
port 710 nsew ground bidirectional
rlabel metal5 s -2936 271876 586860 272476 6 vssd1
port 711 nsew ground bidirectional
rlabel metal5 s -2936 235876 586860 236476 6 vssd1
port 712 nsew ground bidirectional
rlabel metal5 s -2936 199876 586860 200476 6 vssd1
port 713 nsew ground bidirectional
rlabel metal5 s -2936 163876 586860 164476 6 vssd1
port 714 nsew ground bidirectional
rlabel metal5 s -2936 127876 586860 128476 6 vssd1
port 715 nsew ground bidirectional
rlabel metal5 s -2936 91876 586860 92476 6 vssd1
port 716 nsew ground bidirectional
rlabel metal5 s -2936 55876 586860 56476 6 vssd1
port 717 nsew ground bidirectional
rlabel metal5 s -2936 19876 586860 20476 6 vssd1
port 718 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 719 nsew ground bidirectional
rlabel metal4 s 580404 -3744 581004 707680 6 vccd2
port 720 nsew power bidirectional
rlabel metal4 s 544404 -3744 545004 707680 6 vccd2
port 721 nsew power bidirectional
rlabel metal4 s 508404 -3744 509004 707680 6 vccd2
port 722 nsew power bidirectional
rlabel metal4 s 472404 -3744 473004 707680 6 vccd2
port 723 nsew power bidirectional
rlabel metal4 s 436404 -3744 437004 707680 6 vccd2
port 724 nsew power bidirectional
rlabel metal4 s 400404 -3744 401004 707680 6 vccd2
port 725 nsew power bidirectional
rlabel metal4 s 364404 -3744 365004 707680 6 vccd2
port 726 nsew power bidirectional
rlabel metal4 s 328404 -3744 329004 707680 6 vccd2
port 727 nsew power bidirectional
rlabel metal4 s 292404 421000 293004 707680 6 vccd2
port 728 nsew power bidirectional
rlabel metal4 s 256404 421000 257004 707680 6 vccd2
port 729 nsew power bidirectional
rlabel metal4 s 220404 -3744 221004 707680 6 vccd2
port 730 nsew power bidirectional
rlabel metal4 s 184404 -3744 185004 707680 6 vccd2
port 731 nsew power bidirectional
rlabel metal4 s 148404 -3744 149004 707680 6 vccd2
port 732 nsew power bidirectional
rlabel metal4 s 112404 -3744 113004 707680 6 vccd2
port 733 nsew power bidirectional
rlabel metal4 s 76404 -3744 77004 707680 6 vccd2
port 734 nsew power bidirectional
rlabel metal4 s 40404 -3744 41004 707680 6 vccd2
port 735 nsew power bidirectional
rlabel metal4 s 4404 -3744 5004 707680 6 vccd2
port 736 nsew power bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 737 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 738 nsew power bidirectional
rlabel metal4 s 292404 -3744 293004 329000 6 vccd2
port 739 nsew power bidirectional
rlabel metal4 s 256404 -3744 257004 329000 6 vccd2
port 740 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2
port 741 nsew power bidirectional
rlabel metal5 s -4816 689476 588740 690076 6 vccd2
port 742 nsew power bidirectional
rlabel metal5 s -4816 653476 588740 654076 6 vccd2
port 743 nsew power bidirectional
rlabel metal5 s -4816 617476 588740 618076 6 vccd2
port 744 nsew power bidirectional
rlabel metal5 s -4816 581476 588740 582076 6 vccd2
port 745 nsew power bidirectional
rlabel metal5 s -4816 545476 588740 546076 6 vccd2
port 746 nsew power bidirectional
rlabel metal5 s -4816 509476 588740 510076 6 vccd2
port 747 nsew power bidirectional
rlabel metal5 s -4816 473476 588740 474076 6 vccd2
port 748 nsew power bidirectional
rlabel metal5 s -4816 437476 588740 438076 6 vccd2
port 749 nsew power bidirectional
rlabel metal5 s -4816 401476 588740 402076 6 vccd2
port 750 nsew power bidirectional
rlabel metal5 s -4816 365476 588740 366076 6 vccd2
port 751 nsew power bidirectional
rlabel metal5 s -4816 329476 588740 330076 6 vccd2
port 752 nsew power bidirectional
rlabel metal5 s -4816 293476 588740 294076 6 vccd2
port 753 nsew power bidirectional
rlabel metal5 s -4816 257476 588740 258076 6 vccd2
port 754 nsew power bidirectional
rlabel metal5 s -4816 221476 588740 222076 6 vccd2
port 755 nsew power bidirectional
rlabel metal5 s -4816 185476 588740 186076 6 vccd2
port 756 nsew power bidirectional
rlabel metal5 s -4816 149476 588740 150076 6 vccd2
port 757 nsew power bidirectional
rlabel metal5 s -4816 113476 588740 114076 6 vccd2
port 758 nsew power bidirectional
rlabel metal5 s -4816 77476 588740 78076 6 vccd2
port 759 nsew power bidirectional
rlabel metal5 s -4816 41476 588740 42076 6 vccd2
port 760 nsew power bidirectional
rlabel metal5 s -4816 5476 588740 6076 6 vccd2
port 761 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 762 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 763 nsew ground bidirectional
rlabel metal4 s 562404 -3744 563004 707680 6 vssd2
port 764 nsew ground bidirectional
rlabel metal4 s 526404 -3744 527004 707680 6 vssd2
port 765 nsew ground bidirectional
rlabel metal4 s 490404 -3744 491004 707680 6 vssd2
port 766 nsew ground bidirectional
rlabel metal4 s 454404 -3744 455004 707680 6 vssd2
port 767 nsew ground bidirectional
rlabel metal4 s 418404 -3744 419004 707680 6 vssd2
port 768 nsew ground bidirectional
rlabel metal4 s 382404 -3744 383004 707680 6 vssd2
port 769 nsew ground bidirectional
rlabel metal4 s 346404 -3744 347004 707680 6 vssd2
port 770 nsew ground bidirectional
rlabel metal4 s 310404 421000 311004 707680 6 vssd2
port 771 nsew ground bidirectional
rlabel metal4 s 274404 421000 275004 707680 6 vssd2
port 772 nsew ground bidirectional
rlabel metal4 s 238404 421000 239004 707680 6 vssd2
port 773 nsew ground bidirectional
rlabel metal4 s 202404 -3744 203004 707680 6 vssd2
port 774 nsew ground bidirectional
rlabel metal4 s 166404 -3744 167004 707680 6 vssd2
port 775 nsew ground bidirectional
rlabel metal4 s 130404 -3744 131004 707680 6 vssd2
port 776 nsew ground bidirectional
rlabel metal4 s 94404 -3744 95004 707680 6 vssd2
port 777 nsew ground bidirectional
rlabel metal4 s 58404 -3744 59004 707680 6 vssd2
port 778 nsew ground bidirectional
rlabel metal4 s 22404 -3744 23004 707680 6 vssd2
port 779 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 780 nsew ground bidirectional
rlabel metal4 s 310404 -3744 311004 329000 6 vssd2
port 781 nsew ground bidirectional
rlabel metal4 s 274404 -3744 275004 329000 6 vssd2
port 782 nsew ground bidirectional
rlabel metal4 s 238404 -3744 239004 329000 6 vssd2
port 783 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2
port 784 nsew ground bidirectional
rlabel metal5 s -4816 671476 588740 672076 6 vssd2
port 785 nsew ground bidirectional
rlabel metal5 s -4816 635476 588740 636076 6 vssd2
port 786 nsew ground bidirectional
rlabel metal5 s -4816 599476 588740 600076 6 vssd2
port 787 nsew ground bidirectional
rlabel metal5 s -4816 563476 588740 564076 6 vssd2
port 788 nsew ground bidirectional
rlabel metal5 s -4816 527476 588740 528076 6 vssd2
port 789 nsew ground bidirectional
rlabel metal5 s -4816 491476 588740 492076 6 vssd2
port 790 nsew ground bidirectional
rlabel metal5 s -4816 455476 588740 456076 6 vssd2
port 791 nsew ground bidirectional
rlabel metal5 s -4816 419476 588740 420076 6 vssd2
port 792 nsew ground bidirectional
rlabel metal5 s -4816 383476 588740 384076 6 vssd2
port 793 nsew ground bidirectional
rlabel metal5 s -4816 347476 588740 348076 6 vssd2
port 794 nsew ground bidirectional
rlabel metal5 s -4816 311476 588740 312076 6 vssd2
port 795 nsew ground bidirectional
rlabel metal5 s -4816 275476 588740 276076 6 vssd2
port 796 nsew ground bidirectional
rlabel metal5 s -4816 239476 588740 240076 6 vssd2
port 797 nsew ground bidirectional
rlabel metal5 s -4816 203476 588740 204076 6 vssd2
port 798 nsew ground bidirectional
rlabel metal5 s -4816 167476 588740 168076 6 vssd2
port 799 nsew ground bidirectional
rlabel metal5 s -4816 131476 588740 132076 6 vssd2
port 800 nsew ground bidirectional
rlabel metal5 s -4816 95476 588740 96076 6 vssd2
port 801 nsew ground bidirectional
rlabel metal5 s -4816 59476 588740 60076 6 vssd2
port 802 nsew ground bidirectional
rlabel metal5 s -4816 23476 588740 24076 6 vssd2
port 803 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 804 nsew ground bidirectional
rlabel metal4 s 548004 -5624 548604 709560 6 vdda1
port 805 nsew power bidirectional
rlabel metal4 s 512004 -5624 512604 709560 6 vdda1
port 806 nsew power bidirectional
rlabel metal4 s 476004 -5624 476604 709560 6 vdda1
port 807 nsew power bidirectional
rlabel metal4 s 440004 -5624 440604 709560 6 vdda1
port 808 nsew power bidirectional
rlabel metal4 s 404004 -5624 404604 709560 6 vdda1
port 809 nsew power bidirectional
rlabel metal4 s 368004 -5624 368604 709560 6 vdda1
port 810 nsew power bidirectional
rlabel metal4 s 332004 -5624 332604 709560 6 vdda1
port 811 nsew power bidirectional
rlabel metal4 s 296004 421000 296604 709560 6 vdda1
port 812 nsew power bidirectional
rlabel metal4 s 260004 421000 260604 709560 6 vdda1
port 813 nsew power bidirectional
rlabel metal4 s 224004 -5624 224604 709560 6 vdda1
port 814 nsew power bidirectional
rlabel metal4 s 188004 -5624 188604 709560 6 vdda1
port 815 nsew power bidirectional
rlabel metal4 s 152004 -5624 152604 709560 6 vdda1
port 816 nsew power bidirectional
rlabel metal4 s 116004 -5624 116604 709560 6 vdda1
port 817 nsew power bidirectional
rlabel metal4 s 80004 -5624 80604 709560 6 vdda1
port 818 nsew power bidirectional
rlabel metal4 s 44004 -5624 44604 709560 6 vdda1
port 819 nsew power bidirectional
rlabel metal4 s 8004 -5624 8604 709560 6 vdda1
port 820 nsew power bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 821 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 822 nsew power bidirectional
rlabel metal4 s 296004 -5624 296604 329000 6 vdda1
port 823 nsew power bidirectional
rlabel metal4 s 260004 -5624 260604 329000 6 vdda1
port 824 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1
port 825 nsew power bidirectional
rlabel metal5 s -6696 693076 590620 693676 6 vdda1
port 826 nsew power bidirectional
rlabel metal5 s -6696 657076 590620 657676 6 vdda1
port 827 nsew power bidirectional
rlabel metal5 s -6696 621076 590620 621676 6 vdda1
port 828 nsew power bidirectional
rlabel metal5 s -6696 585076 590620 585676 6 vdda1
port 829 nsew power bidirectional
rlabel metal5 s -6696 549076 590620 549676 6 vdda1
port 830 nsew power bidirectional
rlabel metal5 s -6696 513076 590620 513676 6 vdda1
port 831 nsew power bidirectional
rlabel metal5 s -6696 477076 590620 477676 6 vdda1
port 832 nsew power bidirectional
rlabel metal5 s -6696 441076 590620 441676 6 vdda1
port 833 nsew power bidirectional
rlabel metal5 s -6696 405076 590620 405676 6 vdda1
port 834 nsew power bidirectional
rlabel metal5 s -6696 369076 590620 369676 6 vdda1
port 835 nsew power bidirectional
rlabel metal5 s -6696 333076 590620 333676 6 vdda1
port 836 nsew power bidirectional
rlabel metal5 s -6696 297076 590620 297676 6 vdda1
port 837 nsew power bidirectional
rlabel metal5 s -6696 261076 590620 261676 6 vdda1
port 838 nsew power bidirectional
rlabel metal5 s -6696 225076 590620 225676 6 vdda1
port 839 nsew power bidirectional
rlabel metal5 s -6696 189076 590620 189676 6 vdda1
port 840 nsew power bidirectional
rlabel metal5 s -6696 153076 590620 153676 6 vdda1
port 841 nsew power bidirectional
rlabel metal5 s -6696 117076 590620 117676 6 vdda1
port 842 nsew power bidirectional
rlabel metal5 s -6696 81076 590620 81676 6 vdda1
port 843 nsew power bidirectional
rlabel metal5 s -6696 45076 590620 45676 6 vdda1
port 844 nsew power bidirectional
rlabel metal5 s -6696 9076 590620 9676 6 vdda1
port 845 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 846 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 847 nsew ground bidirectional
rlabel metal4 s 566004 -5624 566604 709560 6 vssa1
port 848 nsew ground bidirectional
rlabel metal4 s 530004 -5624 530604 709560 6 vssa1
port 849 nsew ground bidirectional
rlabel metal4 s 494004 -5624 494604 709560 6 vssa1
port 850 nsew ground bidirectional
rlabel metal4 s 458004 -5624 458604 709560 6 vssa1
port 851 nsew ground bidirectional
rlabel metal4 s 422004 -5624 422604 709560 6 vssa1
port 852 nsew ground bidirectional
rlabel metal4 s 386004 -5624 386604 709560 6 vssa1
port 853 nsew ground bidirectional
rlabel metal4 s 350004 -5624 350604 709560 6 vssa1
port 854 nsew ground bidirectional
rlabel metal4 s 314004 421000 314604 709560 6 vssa1
port 855 nsew ground bidirectional
rlabel metal4 s 278004 421000 278604 709560 6 vssa1
port 856 nsew ground bidirectional
rlabel metal4 s 242004 421000 242604 709560 6 vssa1
port 857 nsew ground bidirectional
rlabel metal4 s 206004 -5624 206604 709560 6 vssa1
port 858 nsew ground bidirectional
rlabel metal4 s 170004 -5624 170604 709560 6 vssa1
port 859 nsew ground bidirectional
rlabel metal4 s 134004 -5624 134604 709560 6 vssa1
port 860 nsew ground bidirectional
rlabel metal4 s 98004 -5624 98604 709560 6 vssa1
port 861 nsew ground bidirectional
rlabel metal4 s 62004 -5624 62604 709560 6 vssa1
port 862 nsew ground bidirectional
rlabel metal4 s 26004 -5624 26604 709560 6 vssa1
port 863 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 864 nsew ground bidirectional
rlabel metal4 s 314004 -5624 314604 329000 6 vssa1
port 865 nsew ground bidirectional
rlabel metal4 s 278004 -5624 278604 329000 6 vssa1
port 866 nsew ground bidirectional
rlabel metal4 s 242004 -5624 242604 329000 6 vssa1
port 867 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1
port 868 nsew ground bidirectional
rlabel metal5 s -6696 675076 590620 675676 6 vssa1
port 869 nsew ground bidirectional
rlabel metal5 s -6696 639076 590620 639676 6 vssa1
port 870 nsew ground bidirectional
rlabel metal5 s -6696 603076 590620 603676 6 vssa1
port 871 nsew ground bidirectional
rlabel metal5 s -6696 567076 590620 567676 6 vssa1
port 872 nsew ground bidirectional
rlabel metal5 s -6696 531076 590620 531676 6 vssa1
port 873 nsew ground bidirectional
rlabel metal5 s -6696 495076 590620 495676 6 vssa1
port 874 nsew ground bidirectional
rlabel metal5 s -6696 459076 590620 459676 6 vssa1
port 875 nsew ground bidirectional
rlabel metal5 s -6696 423076 590620 423676 6 vssa1
port 876 nsew ground bidirectional
rlabel metal5 s -6696 387076 590620 387676 6 vssa1
port 877 nsew ground bidirectional
rlabel metal5 s -6696 351076 590620 351676 6 vssa1
port 878 nsew ground bidirectional
rlabel metal5 s -6696 315076 590620 315676 6 vssa1
port 879 nsew ground bidirectional
rlabel metal5 s -6696 279076 590620 279676 6 vssa1
port 880 nsew ground bidirectional
rlabel metal5 s -6696 243076 590620 243676 6 vssa1
port 881 nsew ground bidirectional
rlabel metal5 s -6696 207076 590620 207676 6 vssa1
port 882 nsew ground bidirectional
rlabel metal5 s -6696 171076 590620 171676 6 vssa1
port 883 nsew ground bidirectional
rlabel metal5 s -6696 135076 590620 135676 6 vssa1
port 884 nsew ground bidirectional
rlabel metal5 s -6696 99076 590620 99676 6 vssa1
port 885 nsew ground bidirectional
rlabel metal5 s -6696 63076 590620 63676 6 vssa1
port 886 nsew ground bidirectional
rlabel metal5 s -6696 27076 590620 27676 6 vssa1
port 887 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 888 nsew ground bidirectional
rlabel metal4 s 551604 -7504 552204 711440 6 vdda2
port 889 nsew power bidirectional
rlabel metal4 s 515604 -7504 516204 711440 6 vdda2
port 890 nsew power bidirectional
rlabel metal4 s 479604 -7504 480204 711440 6 vdda2
port 891 nsew power bidirectional
rlabel metal4 s 443604 -7504 444204 711440 6 vdda2
port 892 nsew power bidirectional
rlabel metal4 s 407604 -7504 408204 711440 6 vdda2
port 893 nsew power bidirectional
rlabel metal4 s 371604 -7504 372204 711440 6 vdda2
port 894 nsew power bidirectional
rlabel metal4 s 335604 -7504 336204 711440 6 vdda2
port 895 nsew power bidirectional
rlabel metal4 s 299604 421000 300204 711440 6 vdda2
port 896 nsew power bidirectional
rlabel metal4 s 263604 421000 264204 711440 6 vdda2
port 897 nsew power bidirectional
rlabel metal4 s 227604 -7504 228204 711440 6 vdda2
port 898 nsew power bidirectional
rlabel metal4 s 191604 -7504 192204 711440 6 vdda2
port 899 nsew power bidirectional
rlabel metal4 s 155604 -7504 156204 711440 6 vdda2
port 900 nsew power bidirectional
rlabel metal4 s 119604 -7504 120204 711440 6 vdda2
port 901 nsew power bidirectional
rlabel metal4 s 83604 -7504 84204 711440 6 vdda2
port 902 nsew power bidirectional
rlabel metal4 s 47604 -7504 48204 711440 6 vdda2
port 903 nsew power bidirectional
rlabel metal4 s 11604 -7504 12204 711440 6 vdda2
port 904 nsew power bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 905 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 906 nsew power bidirectional
rlabel metal4 s 299604 -7504 300204 329000 6 vdda2
port 907 nsew power bidirectional
rlabel metal4 s 263604 -7504 264204 329000 6 vdda2
port 908 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2
port 909 nsew power bidirectional
rlabel metal5 s -8576 696676 592500 697276 6 vdda2
port 910 nsew power bidirectional
rlabel metal5 s -8576 660676 592500 661276 6 vdda2
port 911 nsew power bidirectional
rlabel metal5 s -8576 624676 592500 625276 6 vdda2
port 912 nsew power bidirectional
rlabel metal5 s -8576 588676 592500 589276 6 vdda2
port 913 nsew power bidirectional
rlabel metal5 s -8576 552676 592500 553276 6 vdda2
port 914 nsew power bidirectional
rlabel metal5 s -8576 516676 592500 517276 6 vdda2
port 915 nsew power bidirectional
rlabel metal5 s -8576 480676 592500 481276 6 vdda2
port 916 nsew power bidirectional
rlabel metal5 s -8576 444676 592500 445276 6 vdda2
port 917 nsew power bidirectional
rlabel metal5 s -8576 408676 592500 409276 6 vdda2
port 918 nsew power bidirectional
rlabel metal5 s -8576 372676 592500 373276 6 vdda2
port 919 nsew power bidirectional
rlabel metal5 s -8576 336676 592500 337276 6 vdda2
port 920 nsew power bidirectional
rlabel metal5 s -8576 300676 592500 301276 6 vdda2
port 921 nsew power bidirectional
rlabel metal5 s -8576 264676 592500 265276 6 vdda2
port 922 nsew power bidirectional
rlabel metal5 s -8576 228676 592500 229276 6 vdda2
port 923 nsew power bidirectional
rlabel metal5 s -8576 192676 592500 193276 6 vdda2
port 924 nsew power bidirectional
rlabel metal5 s -8576 156676 592500 157276 6 vdda2
port 925 nsew power bidirectional
rlabel metal5 s -8576 120676 592500 121276 6 vdda2
port 926 nsew power bidirectional
rlabel metal5 s -8576 84676 592500 85276 6 vdda2
port 927 nsew power bidirectional
rlabel metal5 s -8576 48676 592500 49276 6 vdda2
port 928 nsew power bidirectional
rlabel metal5 s -8576 12676 592500 13276 6 vdda2
port 929 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 930 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 569604 -7504 570204 711440 6 vssa2
port 932 nsew ground bidirectional
rlabel metal4 s 533604 -7504 534204 711440 6 vssa2
port 933 nsew ground bidirectional
rlabel metal4 s 497604 -7504 498204 711440 6 vssa2
port 934 nsew ground bidirectional
rlabel metal4 s 461604 -7504 462204 711440 6 vssa2
port 935 nsew ground bidirectional
rlabel metal4 s 425604 -7504 426204 711440 6 vssa2
port 936 nsew ground bidirectional
rlabel metal4 s 389604 -7504 390204 711440 6 vssa2
port 937 nsew ground bidirectional
rlabel metal4 s 353604 -7504 354204 711440 6 vssa2
port 938 nsew ground bidirectional
rlabel metal4 s 317604 421000 318204 711440 6 vssa2
port 939 nsew ground bidirectional
rlabel metal4 s 281604 421000 282204 711440 6 vssa2
port 940 nsew ground bidirectional
rlabel metal4 s 245604 421000 246204 711440 6 vssa2
port 941 nsew ground bidirectional
rlabel metal4 s 209604 -7504 210204 711440 6 vssa2
port 942 nsew ground bidirectional
rlabel metal4 s 173604 -7504 174204 711440 6 vssa2
port 943 nsew ground bidirectional
rlabel metal4 s 137604 -7504 138204 711440 6 vssa2
port 944 nsew ground bidirectional
rlabel metal4 s 101604 -7504 102204 711440 6 vssa2
port 945 nsew ground bidirectional
rlabel metal4 s 65604 -7504 66204 711440 6 vssa2
port 946 nsew ground bidirectional
rlabel metal4 s 29604 -7504 30204 711440 6 vssa2
port 947 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 948 nsew ground bidirectional
rlabel metal4 s 317604 -7504 318204 329000 6 vssa2
port 949 nsew ground bidirectional
rlabel metal4 s 281604 -7504 282204 329000 6 vssa2
port 950 nsew ground bidirectional
rlabel metal4 s 245604 -7504 246204 329000 6 vssa2
port 951 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2
port 952 nsew ground bidirectional
rlabel metal5 s -8576 678676 592500 679276 6 vssa2
port 953 nsew ground bidirectional
rlabel metal5 s -8576 642676 592500 643276 6 vssa2
port 954 nsew ground bidirectional
rlabel metal5 s -8576 606676 592500 607276 6 vssa2
port 955 nsew ground bidirectional
rlabel metal5 s -8576 570676 592500 571276 6 vssa2
port 956 nsew ground bidirectional
rlabel metal5 s -8576 534676 592500 535276 6 vssa2
port 957 nsew ground bidirectional
rlabel metal5 s -8576 498676 592500 499276 6 vssa2
port 958 nsew ground bidirectional
rlabel metal5 s -8576 462676 592500 463276 6 vssa2
port 959 nsew ground bidirectional
rlabel metal5 s -8576 426676 592500 427276 6 vssa2
port 960 nsew ground bidirectional
rlabel metal5 s -8576 390676 592500 391276 6 vssa2
port 961 nsew ground bidirectional
rlabel metal5 s -8576 354676 592500 355276 6 vssa2
port 962 nsew ground bidirectional
rlabel metal5 s -8576 318676 592500 319276 6 vssa2
port 963 nsew ground bidirectional
rlabel metal5 s -8576 282676 592500 283276 6 vssa2
port 964 nsew ground bidirectional
rlabel metal5 s -8576 246676 592500 247276 6 vssa2
port 965 nsew ground bidirectional
rlabel metal5 s -8576 210676 592500 211276 6 vssa2
port 966 nsew ground bidirectional
rlabel metal5 s -8576 174676 592500 175276 6 vssa2
port 967 nsew ground bidirectional
rlabel metal5 s -8576 138676 592500 139276 6 vssa2
port 968 nsew ground bidirectional
rlabel metal5 s -8576 102676 592500 103276 6 vssa2
port 969 nsew ground bidirectional
rlabel metal5 s -8576 66676 592500 67276 6 vssa2
port 970 nsew ground bidirectional
rlabel metal5 s -8576 30676 592500 31276 6 vssa2
port 971 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 972 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
