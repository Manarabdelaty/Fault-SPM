* NGSPICE file created from user_proj_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

.subckt user_proj_top clk done mc[0] mc[10] mc[11] mc[12] mc[13] mc[14] mc[15] mc[16]
+ mc[17] mc[18] mc[19] mc[1] mc[20] mc[21] mc[22] mc[23] mc[24] mc[25] mc[26] mc[27]
+ mc[28] mc[29] mc[2] mc[30] mc[31] mc[3] mc[4] mc[5] mc[6] mc[7] mc[8] mc[9] mp[0]
+ mp[10] mp[11] mp[12] mp[13] mp[14] mp[15] mp[16] mp[17] mp[18] mp[19] mp[1] mp[20]
+ mp[21] mp[22] mp[23] mp[24] mp[25] mp[26] mp[27] mp[28] mp[29] mp[2] mp[30] mp[31]
+ mp[3] mp[4] mp[5] mp[6] mp[7] mp[8] mp[9] prod[0] prod[10] prod[11] prod[12] prod[13]
+ prod[14] prod[15] prod[16] prod[17] prod[18] prod[19] prod[1] prod[20] prod[21]
+ prod[22] prod[23] prod[24] prod[25] prod[26] prod[27] prod[28] prod[29] prod[2]
+ prod[30] prod[31] prod[3] prod[4] prod[5] prod[6] prod[7] prod[8] prod[9] prod_sel
+ rst start tck tdi tdo tdo_paden_o tie[0] tie[100] tie[101] tie[102] tie[103] tie[104]
+ tie[105] tie[106] tie[107] tie[108] tie[109] tie[10] tie[110] tie[111] tie[112]
+ tie[113] tie[114] tie[115] tie[116] tie[117] tie[118] tie[119] tie[11] tie[120]
+ tie[121] tie[122] tie[123] tie[124] tie[125] tie[126] tie[127] tie[128] tie[129]
+ tie[12] tie[130] tie[131] tie[132] tie[133] tie[134] tie[135] tie[136] tie[137]
+ tie[138] tie[139] tie[13] tie[140] tie[141] tie[142] tie[143] tie[144] tie[145]
+ tie[146] tie[147] tie[148] tie[149] tie[14] tie[150] tie[151] tie[152] tie[153]
+ tie[154] tie[155] tie[156] tie[157] tie[158] tie[159] tie[15] tie[160] tie[161]
+ tie[162] tie[163] tie[164] tie[165] tie[166] tie[167] tie[168] tie[169] tie[16]
+ tie[17] tie[18] tie[19] tie[1] tie[20] tie[21] tie[22] tie[23] tie[24] tie[25] tie[26]
+ tie[27] tie[28] tie[29] tie[2] tie[30] tie[31] tie[32] tie[33] tie[34] tie[35] tie[36]
+ tie[37] tie[38] tie[39] tie[3] tie[40] tie[41] tie[42] tie[43] tie[44] tie[45] tie[46]
+ tie[47] tie[48] tie[49] tie[4] tie[50] tie[51] tie[52] tie[53] tie[54] tie[55] tie[56]
+ tie[57] tie[58] tie[59] tie[5] tie[60] tie[61] tie[62] tie[63] tie[64] tie[65] tie[66]
+ tie[67] tie[68] tie[69] tie[6] tie[70] tie[71] tie[72] tie[73] tie[74] tie[75] tie[76]
+ tie[77] tie[78] tie[79] tie[7] tie[80] tie[81] tie[82] tie[83] tie[84] tie[85] tie[86]
+ tie[87] tie[88] tie[89] tie[8] tie[90] tie[91] tie[92] tie[93] tie[94] tie[95] tie[96]
+ tie[97] tie[98] tie[99] tie[9] tms trst VPWR VGND
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1506_ __dut__.__uuf__._1548_/A VGND VGND VPWR VPWR __dut__.__uuf__._1506_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_123_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2740_ __dut__._2894_/CLK __dut__._2740_/D __dut__._2512_/Y VGND VGND VPWR
+ VPWR __dut__._2740_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2671_ clkbuf_5_3_0_tck/X __dut__._2671_/D __dut__._2581_/Y VGND VGND VPWR
+ VPWR __dut__._2671_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1437_ __dut__._2155_/B VGND VGND VPWR VPWR __dut__.__uuf__._1437_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2071__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1622_ __dut__._1658_/A1 tie[38] __dut__._1621_/X VGND VGND VPWR VPWR __dut__._2730_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1368_ __dut__._2183_/B VGND VGND VPWR VPWR __dut__.__uuf__._1368_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1553_ __dut__._1555_/A __dut__._2695_/Q VGND VGND VPWR VPWR __dut__._1553_/X
+ sky130_fd_sc_hd__and2_4
Xclkbuf_4_14_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2426_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1299_ __dut__.__uuf__._1286_/X __dut__.__uuf__._1297_/X __dut__._2207_/B
+ __dut__.__uuf__._1298_/X VGND VGND VPWR VPWR __dut__._2206_/A2 sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_opt_1_tck clkbuf_opt_1_tck/A VGND VGND VPWR VPWR clkbuf_opt_1_tck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_73_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1484_ __dut__._1282_/Y mp[23] __dut__._1483_/X VGND VGND VPWR VPWR __dut__._1484_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_133_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1415__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2105_ __dut__._2105_/A __dut__._2105_/B VGND VGND VPWR VPWR __dut__._2105_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2036_ __dut__._2036_/A1 __dut__._2036_/A2 __dut__._2035_/X VGND VGND VPWR
+ VPWR __dut__._2036_/X sky130_fd_sc_hd__a21o_4
XFILLER_139_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_294_ _312_/CLK _294_/D trst VGND VGND VPWR VPWR _294_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2869_ __dut__._2869_/CLK __dut__._2869_/D __dut__._2383_/Y VGND VGND VPWR
+ VPWR __dut__._2869_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_206_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1995__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2352__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_105_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2340_ __dut__.__uuf__._2348_/CLK __dut__._2184_/X __dut__.__uuf__._1356_/X
+ VGND VGND VPWR VPWR __dut__._2185_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2271_ __dut__.__uuf__._2278_/CLK __dut__._2046_/X __dut__.__uuf__._1605_/X
+ VGND VGND VPWR VPWR __dut__._2047_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_141_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1222_ __dut__.__uuf__._1221_/X __dut__.__uuf__._1218_/X __dut__._2237_/B
+ __dut__._2239_/B __dut__.__uuf__._1215_/X VGND VGND VPWR VPWR __dut__._2236_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1153_ __dut__.__uuf__._1147_/X __dut__.__uuf__._1144_/X __dut__._2283_/B
+ __dut__._2285_/B __dut__.__uuf__._1141_/X VGND VGND VPWR VPWR __dut__._2282_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1084_ __dut__.__uuf__._1114_/A VGND VGND VPWR VPWR __dut__.__uuf__._1084_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_103_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1986_ __dut__.__uuf__._1986_/A VGND VGND VPWR VPWR __dut__._2060_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2723_ clkbuf_5_9_0_tck/X __dut__._2723_/D __dut__._2529_/Y VGND VGND VPWR
+ VPWR __dut__._2723_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_144_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2654_ __dut__._2654_/CLK __dut__._2654_/D __dut__._2598_/Y VGND VGND VPWR
+ VPWR __dut__._2654_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2585_ rst VGND VGND VPWR VPWR __dut__._2585_/Y sky130_fd_sc_hd__inv_2
X__dut__._1605_ __dut__._1793_/A __dut__._2721_/Q VGND VGND VPWR VPWR __dut__._1605_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_94_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1536_ __dut__._1282_/Y mc[7] __dut__._1535_/X VGND VGND VPWR VPWR __dut__._1536_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_19_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1467_ _234_/Y __dut__._2673_/Q VGND VGND VPWR VPWR __dut__._1467_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1464__A2 mp[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1398_ __dut__._1398_/A1 __dut__._1396_/X __dut__._1397_/X VGND VGND VPWR
+ VPWR __dut__._2655_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2225__CLK __dut__.__uuf__._2402_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_12_0_tck clkbuf_3_6_0_tck/X VGND VGND VPWR VPWR clkbuf_5_25_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_42_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2019_ __dut__._2029_/A __dut__._2019_/B VGND VGND VPWR VPWR __dut__._2019_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_139_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_277_ _303_/CLK _277_/D VGND VGND VPWR VPWR _277_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_143_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_156_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_323_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1840_ __dut__.__uuf__._1840_/A VGND VGND VPWR VPWR __dut__.__uuf__._1840_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1771_ __dut__.__uuf__._1771_/A VGND VGND VPWR VPWR __dut__.__uuf__._1988_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2614__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2323_ __dut__.__uuf__._2323_/CLK __dut__._2150_/X __dut__.__uuf__._1441_/X
+ VGND VGND VPWR VPWR __dut__._2151_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_145_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2254_ __dut__.__uuf__._2278_/CLK __dut__._2012_/X __dut__.__uuf__._1627_/X
+ VGND VGND VPWR VPWR __dut__._2013_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2185_ VGND VGND VPWR VPWR __dut__.__uuf__._2185_/HI tie[130] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1205_ __dut__.__uuf__._1192_/X __dut__.__uuf__._1204_/X __dut__._2249_/B
+ __dut__._2251_/B __dut__.__uuf__._1200_/X VGND VGND VPWR VPWR __dut__._2248_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1136_ __dut__.__uuf__._1146_/A VGND VGND VPWR VPWR __dut__.__uuf__._1136_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2248__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_114_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2370_ rst VGND VGND VPWR VPWR __dut__._2370_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1321_ __dut__._1325_/A __dut__._2635_/Q VGND VGND VPWR VPWR __dut__._1321_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1067_ __dut__.__uuf__._1058_/X __dut__.__uuf__._1055_/X __dut__._2341_/B
+ __dut__._2343_/B __dut__.__uuf__._1066_/X VGND VGND VPWR VPWR __dut__._2340_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_130_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_200_ _202_/A VGND VGND VPWR VPWR _200_/X sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1969_ __dut__.__uuf__._1969_/A VGND VGND VPWR VPWR __dut__.__uuf__._1969_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_131_ _311_/Q _230_/A VGND VGND VPWR VPWR _131_/Y sky130_fd_sc_hd__nor2_4
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_tck clkbuf_3_1_0_tck/A VGND VGND VPWR VPWR clkbuf_4_3_0_tck/A sky130_fd_sc_hd__clkbuf_1
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2524__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1060__A __dut__.__uuf__._2054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_90 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1434_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_155_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2706_ clkbuf_5_9_0_tck/X __dut__._2706_/D __dut__._2546_/Y VGND VGND VPWR
+ VPWR __dut__._2706_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2637_ __dut__._2357_/B __dut__._2637_/D __dut__._2615_/Y VGND VGND VPWR
+ VPWR __dut__._2637_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2568_ rst VGND VGND VPWR VPWR __dut__._2568_/Y sky130_fd_sc_hd__inv_2
X__dut__._2499_ rst VGND VGND VPWR VPWR __dut__._2499_/Y sky130_fd_sc_hd__inv_2
X__dut__._1519_ _234_/Y __dut__._2686_/Q VGND VGND VPWR VPWR __dut__._1519_/X sky130_fd_sc_hd__and2_4
XFILLER_19_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1603__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2434__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_273_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1428__A2 mp[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2609__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1823_ __dut__.__uuf__._1823_/A __dut__.__uuf__._1823_/B __dut__.__uuf__._1823_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1824_/A sky130_fd_sc_hd__or3_4
XFILLER_60_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1754_ __dut__.__uuf__._1754_/A VGND VGND VPWR VPWR __dut__.__uuf__._1756_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1685_ __dut__._2319_/B __dut__.__uuf__._1681_/X __dut__._2255_/B
+ __dut__.__uuf__._1682_/X VGND VGND VPWR VPWR prod[12] sky130_fd_sc_hd__o22a_4
XFILLER_146_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1870_ __dut__._1870_/A1 tie[162] __dut__._1869_/X VGND VGND VPWR VPWR __dut__._2854_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1364__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2306_ __dut__.__uuf__._2319_/CLK __dut__._2116_/X __dut__.__uuf__._1516_/X
+ VGND VGND VPWR VPWR __dut__._2117_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2237_ __dut__.__uuf__._2282_/CLK __dut__._1978_/X __dut__.__uuf__._1647_/X
+ VGND VGND VPWR VPWR __dut__._1979_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_0_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2168_ VGND VGND VPWR VPWR __dut__.__uuf__._2168_/HI tie[113] sky130_fd_sc_hd__conb_1
X__dut__._2422_ rst VGND VGND VPWR VPWR __dut__._2422_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2099_ VGND VGND VPWR VPWR __dut__.__uuf__._2099_/HI tie[44] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1119_ __dut__.__uuf__._1118_/X __dut__.__uuf__._1114_/X __dut__._2307_/B
+ __dut__._2309_/B __dut__.__uuf__._1111_/X VGND VGND VPWR VPWR __dut__._2306_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._2353_ __dut__._2355_/A __dut__._2353_/B VGND VGND VPWR VPWR __dut__._2353_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_141_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1304_ __dut__._1282_/Y mc[14] __dut__._1303_/X VGND VGND VPWR VPWR __dut__._1304_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2519__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1423__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2284_ __dut__._2356_/A1 __dut__._2284_/A2 __dut__._2283_/X VGND VGND VPWR
+ VPWR __dut__._2284_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_57_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1999_ __dut__._2213_/A __dut__._1999_/B VGND VGND VPWR VPWR __dut__._1999_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2429__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_119_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1470_ __dut__._1496_/X __dut__.__uuf__._1457_/X __dut__._2141_/B
+ __dut__.__uuf__._1463_/X VGND VGND VPWR VPWR __dut__.__uuf__._1470_/X sky130_fd_sc_hd__o22a_4
XFILLER_143_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2800__CLK clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2022_ __dut__.__uuf__._2022_/A VGND VGND VPWR VPWR __dut__.__uuf__._2022_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_57_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1806_ __dut__._1995_/B __dut__._2001_/B VGND VGND VPWR VPWR __dut__.__uuf__._1807_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1737_ __dut__.__uuf__._1730_/A __dut__.__uuf__._1735_/B __dut__.__uuf__._1723_/X
+ VGND VGND VPWR VPWR __dut__._1966_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_147_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1922_ __dut__._2328_/A1 prod[18] __dut__._1921_/X VGND VGND VPWR VPWR __dut__._2880_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1668_ __dut__.__uuf__._1682_/A VGND VGND VPWR VPWR __dut__.__uuf__._1668_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1853_ __dut__._1853_/A __dut__._2845_/Q VGND VGND VPWR VPWR __dut__._1853_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1888__A2 prod[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1599_ __dut__.__uuf__._1599_/A VGND VGND VPWR VPWR __dut__.__uuf__._1599_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1784_ __dut__._1790_/A1 tie[119] __dut__._1783_/X VGND VGND VPWR VPWR __dut__._2811_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_121_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2405_ rst VGND VGND VPWR VPWR __dut__._2405_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2336_ __dut__._2338_/A1 __dut__._2336_/A2 __dut__._2335_/X VGND VGND VPWR
+ VPWR __dut__._2336_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2267_ __dut__._2267_/A __dut__._2267_/B VGND VGND VPWR VPWR __dut__._2267_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1812__A2 tie[133] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_222 psn_inst_psn_buff_228/A VGND VGND VPWR VPWR __dut__._2275_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_211 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1815_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_200 psn_inst_psn_buff_203/A VGND VGND VPWR VPWR __dut__._2066_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._2198_ __dut__._2200_/A1 __dut__._2198_/A2 __dut__._2197_/X VGND VGND VPWR
+ VPWR __dut__._2198_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_244 psn_inst_psn_buff_246/A VGND VGND VPWR VPWR __dut__._1907_/A
+ sky130_fd_sc_hd__buf_2
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_255 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1707_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_233 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2315_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_277 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1617_/A
+ sky130_fd_sc_hd__buf_2
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_288 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2111_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_266 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1663_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_299 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1461_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_129_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1328__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1500__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2309__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_82_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_236_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1522_ __dut__.__uuf__._1564_/A VGND VGND VPWR VPWR __dut__.__uuf__._1522_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1453_ __dut__.__uuf__._1476_/A VGND VGND VPWR VPWR __dut__.__uuf__._1472_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_144_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2622__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1384_ __dut__.__uuf__._1383_/Y __dut__.__uuf__._1362_/X __dut__.__uuf__._1363_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1384_/X sky130_fd_sc_hd__o21a_4
XFILLER_103_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2005_ __dut__.__uuf__._2005_/A VGND VGND VPWR VPWR __dut__.__uuf__._2007_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_122_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2069__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2121_ __dut__._2149_/A __dut__._2121_/B VGND VGND VPWR VPWR __dut__._2121_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2052_ __dut__._2052_/A1 __dut__._2052_/A2 __dut__._2051_/X VGND VGND VPWR
+ VPWR __dut__._2052_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2846__CLK clkbuf_opt_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1905_ __dut__._1905_/A __dut__._2871_/Q VGND VGND VPWR VPWR __dut__._1905_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2885_ __dut__._2885_/CLK __dut__._2885_/D __dut__._2367_/Y VGND VGND VPWR
+ VPWR __dut__._2885_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2532__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1836_ __dut__._1854_/A1 tie[145] __dut__._1835_/X VGND VGND VPWR VPWR __dut__._2837_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1767_ __dut__._2213_/A __dut__._2802_/Q VGND VGND VPWR VPWR __dut__._1767_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1698_ __dut__._1726_/A1 tie[76] __dut__._1697_/X VGND VGND VPWR VPWR __dut__._2768_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_48_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2319_ __dut__._2319_/A __dut__._2319_/B VGND VGND VPWR VPWR __dut__._2319_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2442__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_186_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2281__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_82_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2617__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1505_ __dut__.__uuf__._1516_/A VGND VGND VPWR VPWR __dut__.__uuf__._1505_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2670_ __dut__._2680_/CLK __dut__._2670_/D __dut__._2582_/Y VGND VGND VPWR
+ VPWR __dut__._2670_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1436_ __dut__.__uuf__._1449_/A VGND VGND VPWR VPWR __dut__.__uuf__._1436_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1712__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1621_ __dut__._1661_/A __dut__._2729_/Q VGND VGND VPWR VPWR __dut__._1621_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1367_ __dut__.__uuf__._1393_/A VGND VGND VPWR VPWR __dut__.__uuf__._1367_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1552_ __dut__._1554_/A1 tie[3] __dut__._1551_/X VGND VGND VPWR VPWR __dut__._2695_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1298_ __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR __dut__.__uuf__._1298_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_133_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1483_ _234_/Y __dut__._2677_/Q VGND VGND VPWR VPWR __dut__._1483_/X sky130_fd_sc_hd__and2_4
Xclkbuf_3_6_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0___dut__.__uuf__.__clk_source__/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2104_ __dut__._2104_/A1 __dut__._2104_/A2 __dut__._2103_/X VGND VGND VPWR
+ VPWR __dut__._2104_/X sky130_fd_sc_hd__a21o_4
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2527__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1431__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2035_ __dut__._2051_/A __dut__._2035_/B VGND VGND VPWR VPWR __dut__._2035_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_293_ _303_/CLK _293_/D trst VGND VGND VPWR VPWR _293_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1998__A __dut__.__uuf__._1998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2868_ __dut__._2869_/CLK __dut__._2868_/D __dut__._2384_/Y VGND VGND VPWR
+ VPWR __dut__._2868_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1819_ __dut__._1853_/A __dut__._2828_/Q VGND VGND VPWR VPWR __dut__._1819_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2799_ _271_/CLK __dut__._2799_/D __dut__._2453_/Y VGND VGND VPWR VPWR __dut__._2799_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_96_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._2437__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_101_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2270_ __dut__.__uuf__._2270_/CLK __dut__._2044_/X __dut__.__uuf__._1607_/X
+ VGND VGND VPWR VPWR __dut__._2045_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1221_ __dut__.__uuf__._1478_/A VGND VGND VPWR VPWR __dut__.__uuf__._1221_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_141_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1152_ __dut__.__uuf__._1161_/A VGND VGND VPWR VPWR __dut__.__uuf__._1152_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2691__CLK clkbuf_5_2_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1083_ __dut__.__uuf__._1086_/A VGND VGND VPWR VPWR __dut__.__uuf__._1083_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1985_ __dut__.__uuf__._1985_/A __dut__.__uuf__._1985_/B __dut__.__uuf__._1985_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1986_/A sky130_fd_sc_hd__or3_4
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__308__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2722_ clkbuf_5_8_0_tck/X __dut__._2722_/D __dut__._2530_/Y VGND VGND VPWR
+ VPWR __dut__._2722_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1419_ __dut__._2163_/B VGND VGND VPWR VPWR __dut__.__uuf__._1419_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_144_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2653_ __dut__._2654_/CLK __dut__._2653_/D __dut__._2599_/Y VGND VGND VPWR
+ VPWR __dut__._2653_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2399_ __dut__.__uuf__._2402_/CLK __dut__._2302_/X __dut__.__uuf__._1123_/X
+ VGND VGND VPWR VPWR __dut__._2303_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1604_ __dut__._1604_/A1 tie[29] __dut__._1603_/X VGND VGND VPWR VPWR __dut__._2721_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2584_ rst VGND VGND VPWR VPWR __dut__._2584_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1535_ _234_/Y __dut__._2690_/Q VGND VGND VPWR VPWR __dut__._1535_/X sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_87_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1466_ __dut__._1466_/A1 __dut__._1464_/X __dut__._1465_/X VGND VGND VPWR
+ VPWR __dut__._2672_/D sky130_fd_sc_hd__a21o_4
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1397_ __dut__._2095_/A __dut__._2654_/Q VGND VGND VPWR VPWR __dut__._1397_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2018_ __dut__._2024_/A1 __dut__._2018_/A2 __dut__._2017_/X VGND VGND VPWR
+ VPWR __dut__._2018_/X sky130_fd_sc_hd__a21o_4
X_276_ _193_/A _276_/D VGND VGND VPWR VPWR _276_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_149_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_316_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1770_ __dut__.__uuf__._1761_/A __dut__.__uuf__._1768_/B __dut__.__uuf__._1723_/X
+ VGND VGND VPWR VPWR __dut__._1978_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_60_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1612__B1 __dut__._1611_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2322_ __dut__.__uuf__._2323_/CLK __dut__._2148_/X __dut__.__uuf__._1445_/X
+ VGND VGND VPWR VPWR __dut__._2149_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2253_ __dut__.__uuf__._2278_/CLK __dut__._2010_/X __dut__.__uuf__._1628_/X
+ VGND VGND VPWR VPWR __dut__._2011_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2184_ VGND VGND VPWR VPWR __dut__.__uuf__._2184_/HI tie[129] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1204_ __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR __dut__.__uuf__._1204_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1135_ __dut__.__uuf__._1149_/A VGND VGND VPWR VPWR __dut__.__uuf__._1146_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1320_ __dut__._1282_/Y mc[18] __dut__._1319_/X VGND VGND VPWR VPWR __dut__._1320_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_114_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1066_ __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR __dut__.__uuf__._1066_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2077__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1968_ __dut__._2055_/B __dut__._2061_/B VGND VGND VPWR VPWR __dut__.__uuf__._1969_/A
+ sky130_fd_sc_hd__and2_4
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_130_ _307_/Q VGND VGND VPWR VPWR _130_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1899_ __dut__.__uuf__._1931_/A __dut__.__uuf__._1899_/B __dut__.__uuf__._1899_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1900_/A sky130_fd_sc_hd__or3_4
XFILLER_139_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_91 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1430_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_80 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2142_/A1 sky130_fd_sc_hd__buf_2
XFILLER_105_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2705_ __dut__._2721_/CLK __dut__._2705_/D __dut__._2547_/Y VGND VGND VPWR
+ VPWR __dut__._2705_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2540__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2636_ __dut__._2357_/B __dut__._2636_/D __dut__._2616_/Y VGND VGND VPWR
+ VPWR __dut__._2636_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2567_ rst VGND VGND VPWR VPWR __dut__._2567_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2498_ rst VGND VGND VPWR VPWR __dut__._2498_/Y sky130_fd_sc_hd__inv_2
X__dut__._1518_ __dut__._1530_/A1 __dut__._1516_/X __dut__._1517_/X VGND VGND VPWR
+ VPWR __dut__._2685_/D sky130_fd_sc_hd__a21o_4
XFILLER_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1449_ __dut__._1449_/A __dut__._2667_/Q VGND VGND VPWR VPWR __dut__._1449_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_259_ _193_/A _259_/D VGND VGND VPWR VPWR _259_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_143_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2450__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_266_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1248__A1 __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1822_ __dut__.__uuf__._1821_/X __dut__.__uuf__._1819_/B __dut__.__uuf__._1819_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1823_/C sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._2625__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1753_ __dut__.__uuf__._1798_/A __dut__.__uuf__._1753_/B __dut__.__uuf__._1753_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1754_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1684_ __dut__._2317_/B __dut__.__uuf__._1681_/X __dut__._2253_/B
+ __dut__.__uuf__._1682_/X VGND VGND VPWR VPWR prod[11] sky130_fd_sc_hd__o22a_4
XFILLER_109_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1364__A2 mc[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2305_ __dut__.__uuf__._2319_/CLK __dut__._2114_/X __dut__.__uuf__._1521_/X
+ VGND VGND VPWR VPWR __dut__._2115_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2360__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2236_ __dut__.__uuf__._2282_/CLK __dut__._1976_/X __dut__.__uuf__._1648_/X
+ VGND VGND VPWR VPWR __dut__._1977_/B sky130_fd_sc_hd__dfrtp_4
Xclkbuf_4_11_0_tck clkbuf_3_5_0_tck/X VGND VGND VPWR VPWR clkbuf_5_23_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2421_ rst VGND VGND VPWR VPWR __dut__._2421_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2167_ VGND VGND VPWR VPWR __dut__.__uuf__._2167_/HI tie[112] sky130_fd_sc_hd__conb_1
XFILLER_88_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2098_ VGND VGND VPWR VPWR __dut__.__uuf__._2098_/HI tie[43] sky130_fd_sc_hd__conb_1
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1118_ __dut__.__uuf__._1177_/A VGND VGND VPWR VPWR __dut__.__uuf__._1118_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2352_ __dut__._2356_/A1 __dut__._2352_/A2 __dut__._2351_/X VGND VGND VPWR
+ VPWR __dut__._2352_/X sky130_fd_sc_hd__a21o_4
X__dut__._1303_ _234_/Y __dut__._2632_/Q VGND VGND VPWR VPWR __dut__._1303_/X sky130_fd_sc_hd__and2_4
XFILLER_28_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2283_ __dut__._2285_/A __dut__._2283_/B VGND VGND VPWR VPWR __dut__._2283_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1049_ __dut__.__uuf__._1057_/A VGND VGND VPWR VPWR __dut__.__uuf__._1049_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1336__A __dut__.__uuf__._1711_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2535__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1998_ __dut__._2000_/A1 __dut__._1998_/A2 __dut__._1997_/X VGND VGND VPWR
+ VPWR __dut__._1998_/X sky130_fd_sc_hd__a21o_4
XFILLER_140_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2304__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2619_ rst VGND VGND VPWR VPWR __dut__._2619_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2445__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2238__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__144__A3 tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2021_ __dut__._2075_/B __dut__._2081_/B VGND VGND VPWR VPWR __dut__.__uuf__._2022_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_97_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_tck clkbuf_3_1_0_tck/A VGND VGND VPWR VPWR clkbuf_4_1_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1156__A __dut__.__uuf__._1215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1805_ __dut__._1540_/X VGND VGND VPWR VPWR __dut__.__uuf__._1809_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_138_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1736_ __dut__.__uuf__._1736_/A VGND VGND VPWR VPWR __dut__._1968_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1921_ __dut__._2327_/A __dut__._2879_/Q VGND VGND VPWR VPWR __dut__._1921_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1667_ __dut__._1528_/X VGND VGND VPWR VPWR __dut__.__uuf__._1682_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1852_ __dut__._1854_/A1 tie[153] __dut__._1851_/X VGND VGND VPWR VPWR __dut__._2845_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1598_ __dut__.__uuf__._1599_/A VGND VGND VPWR VPWR __dut__.__uuf__._1598_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_136_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1783_ __dut__._2213_/A __dut__._2810_/Q VGND VGND VPWR VPWR __dut__._1783_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2219_ VGND VGND VPWR VPWR __dut__.__uuf__._2219_/HI tie[164] sky130_fd_sc_hd__conb_1
XFILLER_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2404_ rst VGND VGND VPWR VPWR __dut__._2404_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2335_ __dut__._2335_/A __dut__._2335_/B VGND VGND VPWR VPWR __dut__._2335_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_90_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1066__A __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2266_ __dut__._2266_/A1 __dut__._2266_/A2 __dut__._2265_/X VGND VGND VPWR
+ VPWR __dut__._2266_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2197_ __dut__._2213_/A __dut__._2197_/B VGND VGND VPWR VPWR __dut__._2197_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_201 psn_inst_psn_buff_203/A VGND VGND VPWR VPWR __dut__._2068_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_212 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1813_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_245 psn_inst_psn_buff_246/A VGND VGND VPWR VPWR __dut__._1733_/A
+ sky130_fd_sc_hd__buf_2
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_234 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2321_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_223 psn_inst_psn_buff_228/A VGND VGND VPWR VPWR __dut__._2277_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_278 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1493_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_289 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2109_/A
+ sky130_fd_sc_hd__buf_2
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_256 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1705_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_267 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1949_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_145_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1328__A2 mc[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1609__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1500__A2 mp[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_131_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_229_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1521_ __dut__.__uuf__._1537_/A VGND VGND VPWR VPWR __dut__.__uuf__._1521_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_156_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2798__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1452_ __dut__.__uuf__._1221_/X __dut__.__uuf__._1450_/X __dut__._2147_/B
+ __dut__.__uuf__._2050_/B __dut__.__uuf__._1451_/X VGND VGND VPWR VPWR __dut__._2146_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_104_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1519__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1383_ __dut__._2177_/B VGND VGND VPWR VPWR __dut__.__uuf__._1383_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_103_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2004_ __dut__.__uuf__._2014_/A __dut__.__uuf__._2004_/B __dut__.__uuf__._2004_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2005_/A sky130_fd_sc_hd__or3_4
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2120_ __dut__._2136_/A1 __dut__._2120_/A2 __dut__._2119_/X VGND VGND VPWR
+ VPWR __dut__._2120_/X sky130_fd_sc_hd__a21o_4
XFILLER_38_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2051_ __dut__._2051_/A __dut__._2051_/B VGND VGND VPWR VPWR __dut__._2051_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2085__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1719_ __dut__.__uuf__._1719_/A VGND VGND VPWR VPWR __dut__.__uuf__._1721_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1904_ __dut__._1904_/A1 prod[9] __dut__._1903_/X VGND VGND VPWR VPWR __dut__._2871_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2884_ __dut__._2892_/CLK __dut__._2884_/D __dut__._2368_/Y VGND VGND VPWR
+ VPWR __dut__._2884_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1835_ __dut__._1853_/A __dut__._2836_/Q VGND VGND VPWR VPWR __dut__._1835_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_147_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1766_ __dut__._1766_/A1 tie[110] __dut__._1765_/X VGND VGND VPWR VPWR __dut__._2802_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1697_ __dut__._1701_/A __dut__._2767_/Q VGND VGND VPWR VPWR __dut__._1697_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_3_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2318_ __dut__._2322_/A1 __dut__._2318_/A2 __dut__._2317_/X VGND VGND VPWR
+ VPWR __dut__._2318_/X sky130_fd_sc_hd__a21o_4
X__dut__._2249_ __dut__._2251_/A __dut__._2249_/B VGND VGND VPWR VPWR __dut__._2249_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1339__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_179_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1504_ __dut__.__uuf__._1501_/X __dut__.__uuf__._1495_/X __dut__._2125_/B
+ __dut__.__uuf__._1484_/X __dut__.__uuf__._1503_/X VGND VGND VPWR VPWR __dut__._2124_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1435_ __dut__.__uuf__._1429_/X __dut__.__uuf__._1434_/X __dut__._2155_/B
+ __dut__.__uuf__._1429_/X VGND VGND VPWR VPWR __dut__._2154_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1620_ __dut__._1658_/A1 tie[37] __dut__._1619_/X VGND VGND VPWR VPWR __dut__._2729_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1366_ __dut__.__uuf__._1375_/A VGND VGND VPWR VPWR __dut__.__uuf__._1366_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1551_ __dut__._1555_/A __dut__._2694_/Q VGND VGND VPWR VPWR __dut__._1551_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_86_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0___dut__.__uuf__.__clk_source___A __dut__._2358_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1297_ __dut__.__uuf__._1296_/Y __dut__.__uuf__._2047_/A __dut__.__uuf__._1283_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1297_/X sky130_fd_sc_hd__o21a_4
XFILLER_133_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1476__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1482_ __dut__._1616_/A1 __dut__._1480_/X __dut__._1481_/X VGND VGND VPWR
+ VPWR __dut__._2676_/D sky130_fd_sc_hd__a21o_4
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2103_ __dut__._2103_/A __dut__._2103_/B VGND VGND VPWR VPWR __dut__._2103_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2034_ __dut__._2036_/A1 __dut__._2034_/A2 __dut__._2033_/X VGND VGND VPWR
+ VPWR __dut__._2034_/X sky130_fd_sc_hd__a21o_4
X_292_ _303_/CLK _292_/D trst VGND VGND VPWR VPWR _292_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_psn_inst_psn_buff_32_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1400__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2543__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2867_ __dut__._2869_/CLK __dut__._2867_/D __dut__._2385_/Y VGND VGND VPWR
+ VPWR __dut__._2867_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1818_ __dut__._1854_/A1 tie[136] __dut__._1817_/X VGND VGND VPWR VPWR __dut__._2828_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2798_ _271_/CLK __dut__._2798_/D __dut__._2454_/Y VGND VGND VPWR VPWR __dut__._2798_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_96_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1749_ __dut__._1853_/A __dut__._2793_/Q VGND VGND VPWR VPWR __dut__._1749_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._2453__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1942__A2 prod[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_296_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1220_ __dut__.__uuf__._1220_/A VGND VGND VPWR VPWR __dut__.__uuf__._1220_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_141_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1151_ __dut__.__uuf__._1147_/X __dut__.__uuf__._1144_/X __dut__._2285_/B
+ __dut__._2287_/B __dut__.__uuf__._1141_/X VGND VGND VPWR VPWR __dut__._2284_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._2836__CLK __dut__._2845_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1082_ __dut__.__uuf__._1072_/X __dut__.__uuf__._1069_/X __dut__._2331_/B
+ __dut__._2333_/B __dut__.__uuf__._1081_/X VGND VGND VPWR VPWR __dut__._2330_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_95_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1164__A __dut__.__uuf__._1655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1984_ __dut__.__uuf__._1983_/X __dut__.__uuf__._1981_/B __dut__.__uuf__._1981_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1985_/C sky130_fd_sc_hd__o21a_4
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2363__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2721_ __dut__._2721_/CLK __dut__._2721_/D __dut__._2531_/Y VGND VGND VPWR
+ VPWR __dut__._2721_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1418_ __dut__.__uuf__._1429_/A VGND VGND VPWR VPWR __dut__.__uuf__._1418_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_120_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2398_ __dut__.__uuf__._2398_/CLK __dut__._2300_/X __dut__.__uuf__._1125_/X
+ VGND VGND VPWR VPWR __dut__._2301_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2652_ __dut__._2654_/CLK __dut__._2652_/D __dut__._2600_/Y VGND VGND VPWR
+ VPWR __dut__._2652_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_144_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1349_ __dut__.__uuf__._1342_/X __dut__.__uuf__._1348_/X __dut__._2189_/B
+ __dut__.__uuf__._1342_/X VGND VGND VPWR VPWR __dut__._2188_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1603_ __dut__._1793_/A __dut__._2720_/Q VGND VGND VPWR VPWR __dut__._1603_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2583_ rst VGND VGND VPWR VPWR __dut__._2583_/Y sky130_fd_sc_hd__inv_2
X__dut__._1534_ __dut__._1534_/A1 __dut__._1532_/X __dut__._1533_/X VGND VGND VPWR
+ VPWR __dut__._2689_/D sky130_fd_sc_hd__a21o_4
XFILLER_100_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1465_ __dut__._1465_/A __dut__._2670_/Q VGND VGND VPWR VPWR __dut__._1465_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_85_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1396_ __dut__._1282_/Y mp[3] __dut__._1395_/X VGND VGND VPWR VPWR __dut__._1396_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2538__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1074__A __dut__.__uuf__._2054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2017_ __dut__._2029_/A __dut__._2017_/B VGND VGND VPWR VPWR __dut__._2017_/X
+ sky130_fd_sc_hd__and2_4
X_275_ _193_/A _275_/D VGND VGND VPWR VPWR _275_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2859__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2448__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_211_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_309_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0___dut__.__uuf__.__clk_source__ clkbuf_4_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2270_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2321_ __dut__.__uuf__._2323_/CLK __dut__._2146_/X __dut__.__uuf__._1449_/X
+ VGND VGND VPWR VPWR __dut__._2147_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2252_ __dut__.__uuf__._2278_/CLK __dut__._2008_/X __dut__.__uuf__._1629_/X
+ VGND VGND VPWR VPWR __dut__._2009_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1203_ __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR __dut__.__uuf__._1495_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2183_ VGND VGND VPWR VPWR __dut__.__uuf__._2183_/HI tie[128] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._1527__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1134_ __dut__.__uuf__._1133_/X __dut__.__uuf__._1130_/X __dut__._2297_/B
+ __dut__._2299_/B __dut__.__uuf__._1126_/X VGND VGND VPWR VPWR __dut__._2296_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1065_ __dut__.__uuf__._1071_/A VGND VGND VPWR VPWR __dut__.__uuf__._1065_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_67_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1967_ __dut__._1344_/X VGND VGND VPWR VPWR __dut__.__uuf__._1971_/B
+ sky130_fd_sc_hd__inv_2
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1898_ __dut__.__uuf__._1875_/X __dut__.__uuf__._1896_/B __dut__.__uuf__._1896_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1899_/C sky130_fd_sc_hd__o21a_4
XANTENNA___dut__.__uuf__._2294__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_139_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_92 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1426_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_81 __dut__._1772_/A1 VGND VGND VPWR VPWR psn_inst_psn_buff_99/A
+ sky130_fd_sc_hd__buf_4
Xpsn_inst_psn_buff_70 psn_inst_psn_buff_73/A VGND VGND VPWR VPWR __dut__._2180_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._2704_ __dut__._2721_/CLK __dut__._2704_/D __dut__._2548_/Y VGND VGND VPWR
+ VPWR __dut__._2704_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1726__B1 __dut__.__uuf__._1998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2635_ __dut__._2357_/B __dut__._2635_/D __dut__._2617_/Y VGND VGND VPWR
+ VPWR __dut__._2635_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2566_ rst VGND VGND VPWR VPWR __dut__._2566_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2497_ rst VGND VGND VPWR VPWR __dut__._2497_/Y sky130_fd_sc_hd__inv_2
X__dut__._1517_ __dut__._1517_/A __dut__._2684_/Q VGND VGND VPWR VPWR __dut__._1517_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1842__A1 __dut__._2176_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1448_ __dut__._1282_/Y mp[15] __dut__._1447_/X VGND VGND VPWR VPWR __dut__._1448_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_62_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1379_ _234_/Y __dut__._2651_/Q VGND VGND VPWR VPWR __dut__._1379_/X sky130_fd_sc_hd__and2_4
XFILLER_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_258_ _193_/A _258_/D VGND VGND VPWR VPWR _258_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_189_ _261_/Q _190_/B VGND VGND VPWR VPWR _260_/D sky130_fd_sc_hd__and2_4
XFILLER_143_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1347__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_161_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_259_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1821_ __dut__.__uuf__._2044_/A VGND VGND VPWR VPWR __dut__.__uuf__._1821_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1752_ __dut__._1975_/B __dut__._1981_/B __dut__.__uuf__._1751_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1753_/C sky130_fd_sc_hd__o21ai_4
XFILLER_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1683_ __dut__._2315_/B __dut__.__uuf__._1681_/X __dut__._2251_/B
+ __dut__.__uuf__._1682_/X VGND VGND VPWR VPWR prod[10] sky130_fd_sc_hd__o22a_4
XFILLER_118_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2304_ __dut__.__uuf__._2319_/CLK __dut__._2112_/X __dut__.__uuf__._1526_/X
+ VGND VGND VPWR VPWR __dut__._2113_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2235_ __dut__.__uuf__._2282_/CLK __dut__._1974_/X __dut__.__uuf__._1650_/X
+ VGND VGND VPWR VPWR __dut__._1975_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2166_ VGND VGND VPWR VPWR __dut__.__uuf__._2166_/HI tie[111] sky130_fd_sc_hd__conb_1
X__dut__._2420_ rst VGND VGND VPWR VPWR __dut__._2420_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1117_ __dut__.__uuf__._1191_/A VGND VGND VPWR VPWR __dut__.__uuf__._1177_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2097_ VGND VGND VPWR VPWR __dut__.__uuf__._2097_/HI tie[42] sky130_fd_sc_hd__conb_1
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2351_ __dut__._2355_/A __dut__._2351_/B VGND VGND VPWR VPWR __dut__._2351_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1824__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1302_ __dut__._1346_/A1 __dut__._1300_/X __dut__._1301_/X VGND VGND VPWR
+ VPWR __dut__._2631_/D sky130_fd_sc_hd__a21o_4
X__dut__._2282_ __dut__._2356_/A1 __dut__._2282_/A2 __dut__._2281_/X VGND VGND VPWR
+ VPWR __dut__._2282_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1048_ __dut__.__uuf__._1034_/X __dut__.__uuf__._1038_/X __dut__._2353_/B
+ __dut__._2355_/B __dut__.__uuf__._1040_/X VGND VGND VPWR VPWR __dut__._2352_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2551__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1997_ __dut__._2213_/A __dut__._1997_/B VGND VGND VPWR VPWR __dut__._1997_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2618_ rst VGND VGND VPWR VPWR __dut__._2618_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2549_ rst VGND VGND VPWR VPWR __dut__._2549_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2461__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2020_ __dut__._1364_/X VGND VGND VPWR VPWR __dut__.__uuf__._2024_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_97_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1805__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__270__CLK _270_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1804_ __dut__.__uuf__._1966_/A VGND VGND VPWR VPWR __dut__.__uuf__._1852_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1735_ __dut__.__uuf__._1768_/A __dut__.__uuf__._1735_/B __dut__.__uuf__._1735_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1736_/A sky130_fd_sc_hd__or3_4
XFILLER_138_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1920_ __dut__._2328_/A1 prod[17] __dut__._1919_/X VGND VGND VPWR VPWR __dut__._2879_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1666_ __dut__.__uuf__._1681_/A VGND VGND VPWR VPWR __dut__.__uuf__._1666_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1851_ __dut__._1853_/A __dut__._2844_/Q VGND VGND VPWR VPWR __dut__._1851_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_147_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2371__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1597_ __dut__.__uuf__._1599_/A VGND VGND VPWR VPWR __dut__.__uuf__._1597_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1782_ __dut__._2176_/A1 tie[118] __dut__._1781_/X VGND VGND VPWR VPWR __dut__._2810_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_136_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2298__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2218_ VGND VGND VPWR VPWR __dut__.__uuf__._2218_/HI tie[163] sky130_fd_sc_hd__conb_1
XFILLER_76_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2403_ rst VGND VGND VPWR VPWR __dut__._2403_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2149_ VGND VGND VPWR VPWR __dut__.__uuf__._2149_/HI tie[94] sky130_fd_sc_hd__conb_1
XFILLER_75_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2334_ __dut__._2338_/A1 __dut__._2334_/A2 __dut__._2333_/X VGND VGND VPWR
+ VPWR __dut__._2334_/X sky130_fd_sc_hd__a21o_4
XFILLER_29_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_62_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2265_ __dut__._2265_/A __dut__._2265_/B VGND VGND VPWR VPWR __dut__._2265_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_202 psn_inst_psn_buff_203/A VGND VGND VPWR VPWR __dut__._2000_/A1
+ sky130_fd_sc_hd__buf_8
XFILLER_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2196_ __dut__._2200_/A1 __dut__._2196_/A2 __dut__._2195_/X VGND VGND VPWR
+ VPWR __dut__._2196_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2546__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_213 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1811_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_246 psn_inst_psn_buff_246/A VGND VGND VPWR VPWR __dut__._2327_/A
+ sky130_fd_sc_hd__buf_8
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_235 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2323_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_224 psn_inst_psn_buff_228/A VGND VGND VPWR VPWR __dut__._2279_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_257 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1703_/A
+ sky130_fd_sc_hd__buf_2
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_279 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1489_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_268 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1643_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2456__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_124_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_10_0_tck clkbuf_3_5_0_tck/X VGND VGND VPWR VPWR clkbuf_5_21_0_tck/A sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1520_ __dut__.__uuf__._1581_/A VGND VGND VPWR VPWR __dut__.__uuf__._1537_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2355__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_135_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2191__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1451_ __dut__._1516_/X __dut__.__uuf__._1998_/A __dut__._2149_/B
+ __dut__.__uuf__._1438_/X VGND VGND VPWR VPWR __dut__.__uuf__._1451_/X sky130_fd_sc_hd__o22a_4
XFILLER_144_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1382_ __dut__.__uuf__._1401_/A VGND VGND VPWR VPWR __dut__.__uuf__._1382_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1535__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2003_ __dut__._2067_/B __dut__._2073_/B __dut__.__uuf__._2002_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._2004_/C sky130_fd_sc_hd__o21ai_4
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2366__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2050_ __dut__._2052_/A1 __dut__._2050_/A2 __dut__._2049_/X VGND VGND VPWR
+ VPWR __dut__._2050_/X sky130_fd_sc_hd__a21o_4
XANTENNA__303__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1718_ __dut__.__uuf__._1742_/A __dut__.__uuf__._1718_/B __dut__.__uuf__._1718_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1719_/A sky130_fd_sc_hd__or3_4
XFILLER_154_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1903_ __dut__._1903_/A __dut__._2870_/Q VGND VGND VPWR VPWR __dut__._1903_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1649_ __dut__.__uuf__._1655_/A VGND VGND VPWR VPWR __dut__.__uuf__._1654_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2883_ __dut__._2892_/CLK __dut__._2883_/D __dut__._2369_/Y VGND VGND VPWR
+ VPWR __dut__._2883_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1834_ __dut__._1854_/A1 tie[144] __dut__._1833_/X VGND VGND VPWR VPWR __dut__._2836_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1765_ __dut__._1853_/A __dut__._2801_/Q VGND VGND VPWR VPWR __dut__._1765_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1696_ __dut__._1726_/A1 tie[75] __dut__._1695_/X VGND VGND VPWR VPWR __dut__._2767_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2228__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_91_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2317_ __dut__._2317_/A __dut__._2317_/B VGND VGND VPWR VPWR __dut__._2317_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2248_ __dut__._2248_/A1 __dut__._2248_/A2 __dut__._2247_/X VGND VGND VPWR
+ VPWR __dut__._2248_/X sky130_fd_sc_hd__a21o_4
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2179_ __dut__._2189_/A __dut__._2179_/B VGND VGND VPWR VPWR __dut__._2179_/X
+ sky130_fd_sc_hd__and2_4
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1355__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_241_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_339_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1450__A __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1503_ __dut__._1468_/X __dut__.__uuf__._1502_/X __dut__._2127_/B
+ __dut__.__uuf__._1485_/X VGND VGND VPWR VPWR __dut__.__uuf__._1503_/X sky130_fd_sc_hd__o22a_4
XFILLER_116_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1434_ __dut__.__uuf__._1433_/Y __dut__.__uuf__._1413_/X __dut__.__uuf__._1414_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1434_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1365_ __dut__.__uuf__._1353_/X __dut__.__uuf__._1364_/X __dut__._2183_/B
+ __dut__.__uuf__._1353_/X VGND VGND VPWR VPWR __dut__._2182_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1550_ __dut__._1554_/A1 tie[2] __dut__._1549_/X VGND VGND VPWR VPWR __dut__._2694_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1296_ __dut__._2209_/B VGND VGND VPWR VPWR __dut__.__uuf__._1296_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_100_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1481_ __dut__._1481_/A __dut__._2675_/Q VGND VGND VPWR VPWR __dut__._1481_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1476__A2 mp[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2102_ __dut__._2102_/A1 __dut__._2102_/A2 __dut__._2101_/X VGND VGND VPWR
+ VPWR __dut__._2102_/X sky130_fd_sc_hd__a21o_4
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2033_ __dut__._2051_/A __dut__._2033_/B VGND VGND VPWR VPWR __dut__._2033_/X
+ sky130_fd_sc_hd__and2_4
X_291_ _303_/CLK _291_/D trst VGND VGND VPWR VPWR _291_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_25_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1400__A2 mp[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2866_ __dut__._2869_/CLK __dut__._2866_/D __dut__._2386_/Y VGND VGND VPWR
+ VPWR __dut__._2866_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1817_ __dut__._1817_/A __dut__._2827_/Q VGND VGND VPWR VPWR __dut__._1817_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_96_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2797_ _270_/CLK __dut__._2797_/D __dut__._2455_/Y VGND VGND VPWR VPWR __dut__._2797_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_122_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1748_ __dut__._1854_/A1 tie[101] __dut__._1747_/X VGND VGND VPWR VPWR __dut__._2793_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2638__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__296__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1679_ __dut__._1701_/A __dut__._2758_/Q VGND VGND VPWR VPWR __dut__._1679_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_191_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_289_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1150_ __dut__.__uuf__._1161_/A VGND VGND VPWR VPWR __dut__.__uuf__._1150_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_141_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1081_ __dut__.__uuf__._1141_/A VGND VGND VPWR VPWR __dut__.__uuf__._1081_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1983_ __dut__.__uuf__._1983_/A VGND VGND VPWR VPWR __dut__.__uuf__._1983_/X
+ sky130_fd_sc_hd__buf_2
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2720_ __dut__._2721_/CLK __dut__._2720_/D __dut__._2532_/Y VGND VGND VPWR
+ VPWR __dut__._2720_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2651_ clkbuf_5_3_0_tck/X __dut__._2651_/D __dut__._2601_/Y VGND VGND VPWR
+ VPWR __dut__._2651_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1417_ __dut__.__uuf__._1426_/A VGND VGND VPWR VPWR __dut__.__uuf__._1417_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1602_ __dut__._1602_/A1 tie[28] __dut__._1601_/X VGND VGND VPWR VPWR __dut__._2720_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2397_ __dut__.__uuf__._2398_/CLK __dut__._2298_/X __dut__.__uuf__._1128_/X
+ VGND VGND VPWR VPWR __dut__._2299_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_144_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2582_ rst VGND VGND VPWR VPWR __dut__._2582_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1348_ __dut__.__uuf__._1347_/Y __dut__.__uuf__._1336_/X __dut__.__uuf__._1337_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1348_/X sky130_fd_sc_hd__o21a_4
X__dut__._1533_ __dut__._1533_/A __dut__._2682_/Q VGND VGND VPWR VPWR __dut__._1533_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1279_ __dut__.__uuf__._1276_/X __dut__.__uuf__._2050_/B __dut__._2087_/B
+ __dut__.__uuf__._1040_/X VGND VGND VPWR VPWR __dut__._2214_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1464_ __dut__._1282_/Y mp[18] __dut__._1463_/X VGND VGND VPWR VPWR __dut__._1464_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1395_ _234_/Y __dut__._2655_/Q VGND VGND VPWR VPWR __dut__._1395_/X sky130_fd_sc_hd__and2_4
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2016_ __dut__._2016_/A1 __dut__._2016_/A2 __dut__._2015_/X VGND VGND VPWR
+ VPWR __dut__._2016_/X sky130_fd_sc_hd__a21o_4
X_274_ _193_/A _274_/D VGND VGND VPWR VPWR _274_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._2554__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1090__A __dut__.__uuf__._1655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2849_ clkbuf_5_4_0_tck/X __dut__._2849_/D __dut__._2403_/Y VGND VGND VPWR
+ VPWR __dut__._2849_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_204_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2464__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1376__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2803__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2320_ __dut__.__uuf__._2323_/CLK __dut__._2144_/X __dut__.__uuf__._1454_/X
+ VGND VGND VPWR VPWR __dut__._2145_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_114_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2251_ __dut__.__uuf__._2278_/CLK __dut__._2006_/X __dut__.__uuf__._1630_/X
+ VGND VGND VPWR VPWR __dut__._2007_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1202_ __dut__.__uuf__._1206_/A VGND VGND VPWR VPWR __dut__.__uuf__._1202_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_102_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2182_ VGND VGND VPWR VPWR __dut__.__uuf__._2182_/HI tie[127] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1133_ __dut__.__uuf__._1177_/A VGND VGND VPWR VPWR __dut__.__uuf__._1133_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1064_ __dut__.__uuf__._1058_/X __dut__.__uuf__._1055_/X __dut__._2343_/B
+ __dut__._2345_/B __dut__.__uuf__._1051_/X VGND VGND VPWR VPWR __dut__._2342_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1300__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1543__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1966_ __dut__.__uuf__._1966_/A VGND VGND VPWR VPWR __dut__.__uuf__._2014_/A
+ sky130_fd_sc_hd__buf_2
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2374__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1897_ __dut__.__uuf__._1897_/A VGND VGND VPWR VPWR __dut__.__uuf__._1899_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_137_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_71 psn_inst_psn_buff_73/A VGND VGND VPWR VPWR __dut__._2200_/A1
+ sky130_fd_sc_hd__buf_8
X__dut__._2703_ clkbuf_5_8_0_tck/X __dut__._2703_/D __dut__._2549_/Y VGND VGND VPWR
+ VPWR __dut__._2703_/Q sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_82 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1490_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_60 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2204_/A1 sky130_fd_sc_hd__buf_2
XFILLER_151_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_93 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1422_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2634_ __dut__._2357_/B __dut__._2634_/D __dut__._2618_/Y VGND VGND VPWR
+ VPWR __dut__._2634_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_10_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2412_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__._2565_ rst VGND VGND VPWR VPWR __dut__._2565_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_92_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1516_ __dut__._1282_/Y mp[30] __dut__._1515_/X VGND VGND VPWR VPWR __dut__._1516_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._2496_ rst VGND VGND VPWR VPWR __dut__._2496_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2549__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1453__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1447_ _234_/Y __dut__._2668_/Q VGND VGND VPWR VPWR __dut__._1447_/X sky130_fd_sc_hd__and2_4
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1378_ __dut__._1378_/A1 __dut__._1376_/X __dut__._1377_/X VGND VGND VPWR
+ VPWR __dut__._2650_/D sky130_fd_sc_hd__a21o_4
XFILLER_34_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2826__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_257_ _193_/A _257_/D VGND VGND VPWR VPWR _257_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_188_ _262_/Q _190_/B VGND VGND VPWR VPWR _261_/D sky130_fd_sc_hd__and2_4
XFILLER_143_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._2459__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_154_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1363__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_321_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1820_ __dut__.__uuf__._1820_/A VGND VGND VPWR VPWR __dut__.__uuf__._1823_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_33_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1723__A __dut__.__uuf__._1890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1751_ __dut__.__uuf__._1751_/A VGND VGND VPWR VPWR __dut__.__uuf__._1751_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1682_ __dut__.__uuf__._1682_/A VGND VGND VPWR VPWR __dut__.__uuf__._1682_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_119_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2303_ __dut__.__uuf__._2319_/CLK __dut__._2110_/X __dut__.__uuf__._1531_/X
+ VGND VGND VPWR VPWR __dut__._2111_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2234_ __dut__.__uuf__._2282_/CLK __dut__._1972_/X __dut__.__uuf__._1651_/X
+ VGND VGND VPWR VPWR __dut__._1973_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2165_ VGND VGND VPWR VPWR __dut__.__uuf__._2165_/HI tie[110] sky130_fd_sc_hd__conb_1
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1116_ __dut__.__uuf__._1116_/A VGND VGND VPWR VPWR __dut__.__uuf__._1116_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2369__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2096_ VGND VGND VPWR VPWR __dut__.__uuf__._2096_/HI tie[41] sky130_fd_sc_hd__conb_1
X__dut__._2350_ __dut__._2356_/A1 __dut__._2350_/A2 __dut__._2349_/X VGND VGND VPWR
+ VPWR __dut__._2350_/X sky130_fd_sc_hd__a21o_4
XFILLER_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1301_ __dut__._1301_/A __dut__._2630_/Q VGND VGND VPWR VPWR __dut__._1301_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2281_ __dut__._2349_/A __dut__._2281_/B VGND VGND VPWR VPWR __dut__._2281_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1047_ __dut__.__uuf__._1057_/A VGND VGND VPWR VPWR __dut__.__uuf__._1047_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_71_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2849__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1949_ __dut__._2047_/B __dut__._2053_/B __dut__.__uuf__._1948_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1950_/C sky130_fd_sc_hd__o21ai_4
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1996_ __dut__._2000_/A1 __dut__._1996_/A2 __dut__._1995_/X VGND VGND VPWR
+ VPWR __dut__._1996_/X sky130_fd_sc_hd__a21o_4
XFILLER_125_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1760__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2617_ rst VGND VGND VPWR VPWR __dut__._2617_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1512__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2548_ rst VGND VGND VPWR VPWR __dut__._2548_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_5_31_0_tck clkbuf_5_31_0_tck/A VGND VGND VPWR VPWR __dut__._2845_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2479_ rst VGND VGND VPWR VPWR __dut__._2479_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1911__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1543__A __dut__.__uuf__._1564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_309_ _193_/A _309_/D trst VGND VGND VPWR VPWR _309_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_271_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2284__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1821__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1803_ __dut__.__uuf__._1796_/A __dut__.__uuf__._1801_/B __dut__.__uuf__._1782_/X
+ VGND VGND VPWR VPWR __dut__._1990_/A2 sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1734_ __dut__.__uuf__._1276_/X __dut__.__uuf__._1732_/B __dut__.__uuf__._1732_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1735_/C sky130_fd_sc_hd__o21a_4
XFILLER_138_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1665_ __dut__.__uuf__._1702_/A VGND VGND VPWR VPWR __dut__.__uuf__._1681_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1850_ __dut__._1854_/A1 tie[152] __dut__._1849_/X VGND VGND VPWR VPWR __dut__._2844_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1596_ __dut__.__uuf__._1599_/A VGND VGND VPWR VPWR __dut__.__uuf__._1596_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1781_ __dut__._2213_/A __dut__._2809_/Q VGND VGND VPWR VPWR __dut__._1781_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_136_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1742__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2217_ VGND VGND VPWR VPWR __dut__.__uuf__._2217_/HI tie[162] sky130_fd_sc_hd__conb_1
XFILLER_88_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2402_ rst VGND VGND VPWR VPWR __dut__._2402_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2148_ VGND VGND VPWR VPWR __dut__.__uuf__._2148_/HI tie[93] sky130_fd_sc_hd__conb_1
XFILLER_152_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2079_ VGND VGND VPWR VPWR __dut__.__uuf__._2079_/HI tie[24] sky130_fd_sc_hd__conb_1
X__dut__._2333_ __dut__._2335_/A __dut__._2333_/B VGND VGND VPWR VPWR __dut__._2333_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2671__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2264_ __dut__._2264_/A1 __dut__._2264_/A2 __dut__._2263_/X VGND VGND VPWR
+ VPWR __dut__._2264_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_55_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2195_ __dut__._2213_/A __dut__._2195_/B VGND VGND VPWR VPWR __dut__._2195_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_203 psn_inst_psn_buff_203/A VGND VGND VPWR VPWR __dut__._1980_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_236 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2325_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_225 psn_inst_psn_buff_228/A VGND VGND VPWR VPWR __dut__._2285_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_214 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2341_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_258 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1693_/A
+ sky130_fd_sc_hd__buf_2
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_247 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1905_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_269 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1641_/A
+ sky130_fd_sc_hd__buf_2
Xclkbuf_4_9_0___dut__.__uuf__.__clk_source__ clkbuf_4_9_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2402_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2562__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1979_ __dut__._2213_/A __dut__._1979_/B VGND VGND VPWR VPWR __dut__._1979_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_112_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0___dut__.__uuf__.__clk_source__ clkbuf_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR clkbuf_2_3_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_94_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_psn_inst_psn_buff_117_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2472__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1450_ __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR __dut__.__uuf__._1450_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1724__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1381_ __dut__.__uuf__._1476_/A VGND VGND VPWR VPWR __dut__.__uuf__._1401_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_144_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2694__CLK clkbuf_5_2_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2002_ __dut__.__uuf__._2002_/A VGND VGND VPWR VPWR __dut__.__uuf__._2002_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2382__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1717_ __dut__._1959_/B __dut__._1969_/B __dut__.__uuf__._1716_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1718_/C sky130_fd_sc_hd__o21ai_4
XFILLER_154_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1648_ __dut__.__uuf__._1648_/A VGND VGND VPWR VPWR __dut__.__uuf__._1648_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2882_ __dut__._2892_/CLK __dut__._2882_/D __dut__._2370_/Y VGND VGND VPWR
+ VPWR __dut__._2882_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1902_ __dut__._1902_/A1 prod[8] __dut__._1901_/X VGND VGND VPWR VPWR __dut__._2870_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1833_ __dut__._1853_/A __dut__._2835_/Q VGND VGND VPWR VPWR __dut__._1833_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_107_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1579_ __dut__._1384_/X __dut__.__uuf__._1565_/X __dut__._2089_/B
+ __dut__.__uuf__._1309_/A VGND VGND VPWR VPWR __dut__.__uuf__._1579_/X sky130_fd_sc_hd__o22a_4
X__dut__._1764_ __dut__._1854_/A1 tie[109] __dut__._1763_/X VGND VGND VPWR VPWR __dut__._2801_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1695_ __dut__._1701_/A __dut__._2766_/Q VGND VGND VPWR VPWR __dut__._1695_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_103_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2557__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2316_ __dut__._2322_/A1 __dut__._2316_/A2 __dut__._2315_/X VGND VGND VPWR
+ VPWR __dut__._2316_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2247_ __dut__._2251_/A __dut__._2247_/B VGND VGND VPWR VPWR __dut__._2247_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_32_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2178_ __dut__._2200_/A1 __dut__._2178_/A2 __dut__._2177_/X VGND VGND VPWR
+ VPWR __dut__._2178_/X sky130_fd_sc_hd__a21o_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__.__uuf__._1821__A __dut__.__uuf__._2044_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1706__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2467__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_234_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1371__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2322__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_90_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1502_ __dut__.__uuf__._1565_/A VGND VGND VPWR VPWR __dut__.__uuf__._1502_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1433_ __dut__._2157_/B VGND VGND VPWR VPWR __dut__.__uuf__._1433_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1364_ __dut__.__uuf__._1361_/Y __dut__.__uuf__._1362_/X __dut__.__uuf__._1363_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1364_/X sky130_fd_sc_hd__o21a_4
XFILLER_131_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1295_ __dut__.__uuf__._1295_/A VGND VGND VPWR VPWR __dut__.__uuf__._1295_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1480_ __dut__._1282_/Y mp[22] __dut__._1479_/X VGND VGND VPWR VPWR __dut__._1480_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_85_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2377__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1281__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2101_ __dut__._2101_/A __dut__._2101_/B VGND VGND VPWR VPWR __dut__._2101_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2032_ __dut__._2032_/A1 __dut__._2032_/A2 __dut__._2031_/X VGND VGND VPWR
+ VPWR __dut__._2032_/X sky130_fd_sc_hd__a21o_4
X_290_ _303_/CLK _290_/D trst VGND VGND VPWR VPWR _290_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1048__B2 __dut__.__uuf__._1040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_18_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2865_ __dut__._2865_/CLK __dut__._2865_/D __dut__._2387_/Y VGND VGND VPWR
+ VPWR __dut__._2865_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2796_ _270_/CLK __dut__._2796_/D __dut__._2456_/Y VGND VGND VPWR VPWR __dut__._2796_/Q
+ sky130_fd_sc_hd__dfrtp_4
X__dut__._1816_ __dut__._1854_/A1 tie[135] __dut__._1815_/X VGND VGND VPWR VPWR __dut__._2827_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_123_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1747_ __dut__._1853_/A __dut__._2792_/Q VGND VGND VPWR VPWR __dut__._1747_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1678_ __dut__._1726_/A1 tie[66] __dut__._1677_/X VGND VGND VPWR VPWR __dut__._2758_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2287__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_184_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2352__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1080_ __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR __dut__.__uuf__._1141_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_67_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2197__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1982_ __dut__.__uuf__._1982_/A VGND VGND VPWR VPWR __dut__.__uuf__._1985_/B
+ sky130_fd_sc_hd__inv_2
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2650_ __dut__._2654_/CLK __dut__._2650_/D __dut__._2602_/Y VGND VGND VPWR
+ VPWR __dut__._2650_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2396_ __dut__.__uuf__._2398_/CLK __dut__._2296_/X __dut__.__uuf__._1132_/X
+ VGND VGND VPWR VPWR __dut__._2297_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1416_ __dut__.__uuf__._1404_/X __dut__.__uuf__._1415_/X __dut__._2163_/B
+ __dut__.__uuf__._1404_/X VGND VGND VPWR VPWR __dut__._2162_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2810__D __dut__._2810_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1347_ __dut__._2191_/B VGND VGND VPWR VPWR __dut__.__uuf__._1347_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1601_ __dut__._1793_/A __dut__._2719_/Q VGND VGND VPWR VPWR __dut__._1601_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_120_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2581_ rst VGND VGND VPWR VPWR __dut__._2581_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1532_ __dut__._1282_/Y mc[6] __dut__._1531_/X VGND VGND VPWR VPWR __dut__._1532_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1278_ __dut__.__uuf__._1548_/A VGND VGND VPWR VPWR __dut__.__uuf__._2050_/B
+ sky130_fd_sc_hd__buf_2
XFILLER_74_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1463_ _234_/Y __dut__._2672_/Q VGND VGND VPWR VPWR __dut__._1463_/X sky130_fd_sc_hd__and2_4
XFILLER_100_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1394_ __dut__._1394_/A1 __dut__._1392_/X __dut__._1393_/X VGND VGND VPWR
+ VPWR __dut__._2654_/D sky130_fd_sc_hd__a21o_4
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2015_ __dut__._2029_/A __dut__._2015_/B VGND VGND VPWR VPWR __dut__._2015_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_273_ _288_/CLK _273_/D VGND VGND VPWR VPWR _273_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2570__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2848_ clkbuf_5_4_0_tck/X __dut__._2848_/D __dut__._2404_/Y VGND VGND VPWR
+ VPWR __dut__._2848_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2779_ __dut__._2869_/CLK __dut__._2779_/D __dut__._2473_/Y VGND VGND VPWR
+ VPWR __dut__._2779_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1376__A2 mc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2480__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2250_ __dut__.__uuf__._2288_/CLK __dut__._2004_/X __dut__.__uuf__._1632_/X
+ VGND VGND VPWR VPWR __dut__._2005_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_142_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1201_ __dut__.__uuf__._1192_/X __dut__.__uuf__._1188_/X __dut__._2251_/B
+ __dut__._2253_/B __dut__.__uuf__._1200_/X VGND VGND VPWR VPWR __dut__._2250_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_102_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2181_ VGND VGND VPWR VPWR __dut__.__uuf__._2181_/HI tie[126] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1132_ __dut__.__uuf__._1132_/A VGND VGND VPWR VPWR __dut__.__uuf__._1132_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1063_ __dut__.__uuf__._1071_/A VGND VGND VPWR VPWR __dut__.__uuf__._1063_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_83_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1300__A2 mc[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1965_ __dut__.__uuf__._1958_/A __dut__.__uuf__._1963_/B __dut__.__uuf__._1944_/X
+ VGND VGND VPWR VPWR __dut__._2050_/A2 sky130_fd_sc_hd__o21a_4
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1896_ __dut__.__uuf__._1906_/A __dut__.__uuf__._1896_/B __dut__.__uuf__._1896_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1897_/A sky130_fd_sc_hd__or3_4
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2628__CLK clkbuf_5_2_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2390__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_72 psn_inst_psn_buff_73/A VGND VGND VPWR VPWR __dut__._2176_/A1
+ sky130_fd_sc_hd__buf_8
XFILLER_3_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2702_ __dut__._2721_/CLK __dut__._2702_/D __dut__._2550_/Y VGND VGND VPWR
+ VPWR __dut__._2702_/Q sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_83 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1486_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_50 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2090_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_61 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2206_/A1 sky130_fd_sc_hd__buf_2
XFILLER_151_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_94 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1414_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_132_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2633_ __dut__._2357_/B __dut__._2633_/D __dut__._2619_/Y VGND VGND VPWR
+ VPWR __dut__._2633_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2379_ __dut__.__uuf__._2412_/CLK __dut__._2262_/X __dut__.__uuf__._1182_/X
+ VGND VGND VPWR VPWR __dut__._2263_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_105_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2564_ rst VGND VGND VPWR VPWR __dut__._2564_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_85_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1515_ _234_/Y __dut__._2685_/Q VGND VGND VPWR VPWR __dut__._1515_/X sky130_fd_sc_hd__and2_4
Xclkbuf_3_2_0___dut__.__uuf__.__clk_source__ clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_5_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2495_ rst VGND VGND VPWR VPWR __dut__._2495_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1446_ __dut__._1446_/A1 __dut__._1444_/X __dut__._1445_/X VGND VGND VPWR
+ VPWR __dut__._2667_/D sky130_fd_sc_hd__a21o_4
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1377_ __dut__._2095_/A __dut__._2648_/Q VGND VGND VPWR VPWR __dut__._1377_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2565__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_6_0___dut__.__uuf__.__clk_source___A clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_256_ _308_/CLK _256_/D VGND VGND VPWR VPWR _256_/Q sky130_fd_sc_hd__dfxtp_4
X_187_ _263_/Q _190_/B VGND VGND VPWR VPWR _262_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1909__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1530__A2 __dut__._1528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_147_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_314_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1750_ __dut__._1975_/B __dut__._1981_/B VGND VGND VPWR VPWR __dut__.__uuf__._1751_/A
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2475__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1681_ __dut__.__uuf__._1681_/A VGND VGND VPWR VPWR __dut__.__uuf__._1681_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_146_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1819__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2302_ __dut__.__uuf__._2319_/CLK __dut__._2108_/X __dut__.__uuf__._1534_/X
+ VGND VGND VPWR VPWR __dut__._2109_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2233_ __dut__.__uuf__._2282_/CLK __dut__._1970_/X __dut__.__uuf__._1652_/X
+ VGND VGND VPWR VPWR __dut__._1971_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_130_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._2164_ VGND VGND VPWR VPWR __dut__.__uuf__._2164_/HI tie[109] sky130_fd_sc_hd__conb_1
XFILLER_114_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1115_ __dut__.__uuf__._1103_/X __dut__.__uuf__._1114_/X __dut__._2309_/B
+ __dut__._2311_/B __dut__.__uuf__._1111_/X VGND VGND VPWR VPWR __dut__._2308_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_68_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2095_ VGND VGND VPWR VPWR __dut__.__uuf__._2095_/HI tie[40] sky130_fd_sc_hd__conb_1
X__dut__._1300_ __dut__._1282_/Y mc[13] __dut__._1299_/X VGND VGND VPWR VPWR __dut__._1300_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_83_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2280_ __dut__._2356_/A1 __dut__._2280_/A2 __dut__._2279_/X VGND VGND VPWR
+ VPWR __dut__._2280_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1046_ __dut__.__uuf__._1034_/X __dut__.__uuf__._1038_/X __dut__._2355_/B
+ __dut__._1885_/B __dut__.__uuf__._1040_/X VGND VGND VPWR VPWR __dut__._2354_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_56_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2385__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1948_ __dut__.__uuf__._1948_/A VGND VGND VPWR VPWR __dut__.__uuf__._1948_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1879_ __dut__.__uuf__._1871_/A __dut__.__uuf__._1877_/B __dut__.__uuf__._1836_/X
+ VGND VGND VPWR VPWR __dut__._2018_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1995_ __dut__._2213_/A __dut__._1995_/B VGND VGND VPWR VPWR __dut__._1995_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1512__A2 mp[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2616_ rst VGND VGND VPWR VPWR __dut__._2616_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2547_ rst VGND VGND VPWR VPWR __dut__._2547_/Y sky130_fd_sc_hd__inv_2
X__dut__._2478_ rst VGND VGND VPWR VPWR __dut__._2478_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1429_ __dut__._1433_/A __dut__._2662_/Q VGND VGND VPWR VPWR __dut__._1429_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2295__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_308_ _308_/CLK _308_/D trst VGND VGND VPWR VPWR _308_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_3_5_0_tck_A clkbuf_3_5_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_239_ tms _238_/X _127_/X VGND VGND VPWR VPWR _304_/D sky130_fd_sc_hd__a21o_4
XFILLER_115_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_264_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1802_ __dut__.__uuf__._1802_/A VGND VGND VPWR VPWR __dut__._1992_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_33_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1733_ __dut__.__uuf__._1733_/A VGND VGND VPWR VPWR __dut__.__uuf__._1735_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1664_ __dut__._1528_/X VGND VGND VPWR VPWR __dut__.__uuf__._1702_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1595_ __dut__.__uuf__._1599_/A VGND VGND VPWR VPWR __dut__.__uuf__._1595_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1780_ __dut__._1780_/A1 tie[117] __dut__._1779_/X VGND VGND VPWR VPWR __dut__._2809_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_136_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2216_ VGND VGND VPWR VPWR __dut__.__uuf__._2216_/HI tie[161] sky130_fd_sc_hd__conb_1
XFILLER_88_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2401_ rst VGND VGND VPWR VPWR __dut__._2401_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2147_ VGND VGND VPWR VPWR __dut__.__uuf__._2147_/HI tie[92] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2816__CLK clkbuf_5_0_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2078_ VGND VGND VPWR VPWR __dut__.__uuf__._2078_/HI tie[23] sky130_fd_sc_hd__conb_1
X__dut__._2332_ __dut__._2338_/A1 __dut__._2332_/A2 __dut__._2331_/X VGND VGND VPWR
+ VPWR __dut__._2332_/X sky130_fd_sc_hd__a21o_4
X__dut__._2263_ __dut__._2263_/A __dut__._2263_/B VGND VGND VPWR VPWR __dut__._2263_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1029_ __dut__._2221_/B __dut__.__uuf__._1234_/A __dut__._2217_/B
+ __dut__.__uuf__._1029_/D VGND VGND VPWR VPWR __dut__.__uuf__._2051_/C sky130_fd_sc_hd__or4_4
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_204 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1810_/A1 sky130_fd_sc_hd__buf_2
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2194_ __dut__._2200_/A1 __dut__._2194_/A2 __dut__._2193_/X VGND VGND VPWR
+ VPWR __dut__._2194_/X sky130_fd_sc_hd__a21o_4
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_237 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2265_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA_psn_inst_psn_buff_48_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_226 psn_inst_psn_buff_228/A VGND VGND VPWR VPWR __dut__._2313_/A
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_215 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2339_/A
+ sky130_fd_sc_hd__buf_2
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_259 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1691_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_248 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1903_/A
+ sky130_fd_sc_hd__buf_2
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1459__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1978_ __dut__._1980_/A1 __dut__._1978_/A2 __dut__._1977_/X VGND VGND VPWR
+ VPWR __dut__._1978_/X sky130_fd_sc_hd__a21o_4
XFILLER_3_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1380_ __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR __dut__.__uuf__._1476_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_144_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2839__CLK clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1488__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2001_ __dut__._2067_/B __dut__._2073_/B VGND VGND VPWR VPWR __dut__.__uuf__._2002_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_100_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1412__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1716_ __dut__.__uuf__._1716_/A VGND VGND VPWR VPWR __dut__.__uuf__._1716_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1647_ __dut__.__uuf__._1648_/A VGND VGND VPWR VPWR __dut__.__uuf__._1647_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2881_ __dut__._2892_/CLK __dut__._2881_/D __dut__._2371_/Y VGND VGND VPWR
+ VPWR __dut__._2881_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1901_ __dut__._1901_/A __dut__._2869_/Q VGND VGND VPWR VPWR __dut__._1901_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1832_ __dut__._1854_/A1 tie[143] __dut__._1831_/X VGND VGND VPWR VPWR __dut__._2835_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_135_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_30_0_tck clkbuf_5_31_0_tck/A VGND VGND VPWR VPWR _270_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1578_ __dut__.__uuf__._1578_/A VGND VGND VPWR VPWR __dut__.__uuf__._1890_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_150_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__312__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1763_ __dut__._1853_/A __dut__._2800_/Q VGND VGND VPWR VPWR __dut__._1763_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1694_ __dut__._1694_/A1 tie[74] __dut__._1693_/X VGND VGND VPWR VPWR __dut__._2766_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2315_ __dut__._2315_/A __dut__._2315_/B VGND VGND VPWR VPWR __dut__._2315_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2246_ __dut__._2248_/A1 __dut__._2246_/A2 __dut__._2245_/X VGND VGND VPWR
+ VPWR __dut__._2246_/X sky130_fd_sc_hd__a21o_4
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2177_ __dut__._2189_/A __dut__._2177_/B VGND VGND VPWR VPWR __dut__._2177_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_32_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2573__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1917__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2483__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1501_ __dut__.__uuf__._1564_/A VGND VGND VPWR VPWR __dut__.__uuf__._1501_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_117_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1432_ __dut__.__uuf__._1449_/A VGND VGND VPWR VPWR __dut__.__uuf__._1432_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_2_2_0_tck_A clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1827__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1363_ __dut__.__uuf__._1414_/A VGND VGND VPWR VPWR __dut__.__uuf__._1363_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1294_ __dut__.__uuf__._1286_/X __dut__.__uuf__._1293_/X __dut__._2209_/B
+ __dut__.__uuf__._1286_/X VGND VGND VPWR VPWR __dut__._2208_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2100_ __dut__._2100_/A1 __dut__._2100_/A2 __dut__._2099_/X VGND VGND VPWR
+ VPWR __dut__._2100_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._1194__A __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2031_ __dut__._2031_/A __dut__._2031_/B VGND VGND VPWR VPWR __dut__._2031_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2297__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1048__A2 __dut__.__uuf__._1038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2393__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1936__A2 prod[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2864_ __dut__._2865_/CLK __dut__._2864_/D __dut__._2388_/Y VGND VGND VPWR
+ VPWR __dut__._2864_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2795_ _270_/CLK __dut__._2795_/D __dut__._2457_/Y VGND VGND VPWR VPWR __dut__._2795_/Q
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1737__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1815_ __dut__._1815_/A __dut__._2826_/Q VGND VGND VPWR VPWR __dut__._1815_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_150_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1746_ __dut__._1854_/A1 tie[100] __dut__._1745_/X VGND VGND VPWR VPWR __dut__._2792_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1677_ __dut__._1701_/A __dut__._2757_/Q VGND VGND VPWR VPWR __dut__._1677_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_1_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2568__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2229_ __dut__._2313_/A __dut__._2229_/B VGND VGND VPWR VPWR __dut__._2229_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_177_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2478__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1981_ __dut__.__uuf__._2014_/A __dut__.__uuf__._1981_/B __dut__.__uuf__._1981_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1982_/A sky130_fd_sc_hd__or3_4
XFILLER_149_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2395_ __dut__.__uuf__._2426_/CLK __dut__._2294_/X __dut__.__uuf__._1136_/X
+ VGND VGND VPWR VPWR __dut__._2295_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1415_ __dut__.__uuf__._1412_/Y __dut__.__uuf__._1413_/X __dut__.__uuf__._1414_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1415_/X sky130_fd_sc_hd__o21a_4
XFILLER_132_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1346_ __dut__.__uuf__._1350_/A VGND VGND VPWR VPWR __dut__.__uuf__._1346_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1600_ __dut__._1790_/A1 tie[27] __dut__._1599_/X VGND VGND VPWR VPWR __dut__._2719_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_120_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2580_ rst VGND VGND VPWR VPWR __dut__._2580_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1531_ _234_/Y __dut__._2689_/Q VGND VGND VPWR VPWR __dut__._1531_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1277_ __dut__.__uuf__._1461_/A VGND VGND VPWR VPWR __dut__.__uuf__._1548_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1854__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2388__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1462_ __dut__._1462_/A1 __dut__._1460_/X __dut__._1461_/X VGND VGND VPWR
+ VPWR __dut__._2671_/D sky130_fd_sc_hd__a21o_4
XFILLER_74_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1393_ __dut__._2095_/A __dut__._2653_/Q VGND VGND VPWR VPWR __dut__._1393_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2014_ __dut__._2014_/A1 __dut__._2014_/A2 __dut__._2013_/X VGND VGND VPWR
+ VPWR __dut__._2014_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_0 __dut__._1281_/Y VGND VGND VPWR VPWR __dut__._1772_/A1 sky130_fd_sc_hd__buf_8
XFILLER_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_272_ _288_/CLK _272_/D VGND VGND VPWR VPWR _272_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_psn_inst_psn_buff_30_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2847_ clkbuf_5_4_0_tck/X __dut__._2847_/D __dut__._2405_/Y VGND VGND VPWR
+ VPWR __dut__._2847_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1467__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2312__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2778_ __dut__._2869_/CLK __dut__._2778_/D __dut__._2474_/Y VGND VGND VPWR
+ VPWR __dut__._2778_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_3_1_0___dut__.__uuf__.__clk_source___A clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1729_ __dut__._1729_/A __dut__._2783_/Q VGND VGND VPWR VPWR __dut__._1729_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_294_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1200_ __dut__.__uuf__._1215_/A VGND VGND VPWR VPWR __dut__.__uuf__._1200_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2180_ VGND VGND VPWR VPWR __dut__.__uuf__._2180_/HI tie[125] sky130_fd_sc_hd__conb_1
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1131_ __dut__.__uuf__._1118_/X __dut__.__uuf__._1130_/X __dut__._2299_/B
+ __dut__._2301_/B __dut__.__uuf__._1126_/X VGND VGND VPWR VPWR __dut__._2298_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_102_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1836__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1062_ __dut__.__uuf__._1058_/X __dut__.__uuf__._1055_/X __dut__._2345_/B
+ __dut__._2347_/B __dut__.__uuf__._1051_/X VGND VGND VPWR VPWR __dut__._2344_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_83_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2001__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1964_ __dut__.__uuf__._1964_/A VGND VGND VPWR VPWR __dut__._2052_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1895_ __dut__._2027_/B __dut__._2033_/B __dut__.__uuf__._1894_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1896_/C sky130_fd_sc_hd__o21ai_4
XFILLER_149_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_40 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2058_/A1 sky130_fd_sc_hd__buf_2
XFILLER_152_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1287__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2701_ clkbuf_5_8_0_tck/X __dut__._2701_/D __dut__._2551_/Y VGND VGND VPWR
+ VPWR __dut__._2701_/Q sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_51 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2088_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_73 psn_inst_psn_buff_73/A VGND VGND VPWR VPWR __dut__._2166_/A1
+ sky130_fd_sc_hd__buf_4
Xpsn_inst_psn_buff_62 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2208_/A1 sky130_fd_sc_hd__buf_2
XFILLER_144_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_95 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1410_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_84 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1454_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2378_ __dut__.__uuf__._2412_/CLK __dut__._2260_/X __dut__.__uuf__._1184_/X
+ VGND VGND VPWR VPWR __dut__._2261_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2632_ __dut__._2357_/B __dut__._2632_/D __dut__._2620_/Y VGND VGND VPWR
+ VPWR __dut__._2632_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2563_ rst VGND VGND VPWR VPWR __dut__._2563_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1329_ __dut__.__uuf__._1350_/A VGND VGND VPWR VPWR __dut__.__uuf__._1329_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1514_ __dut__._1530_/A1 __dut__._1512_/X __dut__._1513_/X VGND VGND VPWR
+ VPWR __dut__._2684_/D sky130_fd_sc_hd__a21o_4
XFILLER_101_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2494_ rst VGND VGND VPWR VPWR __dut__._2494_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_78_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1445_ __dut__._1445_/A __dut__._2666_/Q VGND VGND VPWR VPWR __dut__._1445_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_74_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1376_ __dut__._1282_/Y mc[30] __dut__._1375_/X VGND VGND VPWR VPWR __dut__._1376_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_255_ _308_/CLK _255_/D VGND VGND VPWR VPWR _256_/D sky130_fd_sc_hd__dfxtp_4
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2581__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_186_ _264_/Q _186_/B VGND VGND VPWR VPWR _263_/D sky130_fd_sc_hd__or2_4
XFILLER_142_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1925__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_tck_A clkbuf_3_1_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1818__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_307_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1680_ __dut__._2313_/B __dut__.__uuf__._1674_/X __dut__._2249_/B
+ __dut__.__uuf__._1675_/X VGND VGND VPWR VPWR prod[9] sky130_fd_sc_hd__o22a_4
XFILLER_146_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2491__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2301_ __dut__.__uuf__._2319_/CLK __dut__._2106_/X __dut__.__uuf__._1537_/X
+ VGND VGND VPWR VPWR __dut__._2107_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_130_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2232_ __dut__.__uuf__._2348_/CLK __dut__._1968_/X __dut__.__uuf__._1653_/X
+ VGND VGND VPWR VPWR __dut__._1969_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1835__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2163_ VGND VGND VPWR VPWR __dut__.__uuf__._2163_/HI tie[108] sky130_fd_sc_hd__conb_1
XFILLER_87_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2094_ VGND VGND VPWR VPWR __dut__.__uuf__._2094_/HI tie[39] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1114_ __dut__.__uuf__._1114_/A VGND VGND VPWR VPWR __dut__.__uuf__._1114_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_68_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1045_ __dut__.__uuf__._2054_/A VGND VGND VPWR VPWR __dut__.__uuf__._1057_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_83_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2234__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1947_ __dut__._2047_/B __dut__._2053_/B VGND VGND VPWR VPWR __dut__.__uuf__._1948_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1878_ __dut__.__uuf__._1878_/A VGND VGND VPWR VPWR __dut__._2020_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1994_ __dut__._2000_/A1 __dut__._1994_/A2 __dut__._1993_/X VGND VGND VPWR
+ VPWR __dut__._1994_/X sky130_fd_sc_hd__a21o_4
XFILLER_152_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2895__CLK clkbuf_5_0_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2615_ rst VGND VGND VPWR VPWR __dut__._2615_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2546_ rst VGND VGND VPWR VPWR __dut__._2546_/Y sky130_fd_sc_hd__inv_2
X__dut__._2477_ rst VGND VGND VPWR VPWR __dut__._2477_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2576__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1428_ __dut__._1282_/Y mp[10] __dut__._1427_/X VGND VGND VPWR VPWR __dut__._1428_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1359_ _234_/Y __dut__._2646_/Q VGND VGND VPWR VPWR __dut__._1359_/X sky130_fd_sc_hd__and2_4
XFILLER_91_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_307_ _312_/CLK _307_/D trst VGND VGND VPWR VPWR _307_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_238_ _295_/Q _304_/Q VGND VGND VPWR VPWR _238_/X sky130_fd_sc_hd__or2_4
XFILLER_11_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_169_ _278_/Q _171_/B VGND VGND VPWR VPWR _277_/D sky130_fd_sc_hd__or2_4
XFILLER_112_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_257_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2486__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1801_ __dut__.__uuf__._1823_/A __dut__.__uuf__._1801_/B __dut__.__uuf__._1801_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1802_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1732_ __dut__.__uuf__._1742_/A __dut__.__uuf__._1732_/B __dut__.__uuf__._1732_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1733_/A sky130_fd_sc_hd__or3_4
XFILLER_147_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1663_ __dut__.__uuf__._1663_/A VGND VGND VPWR VPWR done sky130_fd_sc_hd__buf_2
XFILLER_146_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1594_ __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR __dut__.__uuf__._1599_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2215_ VGND VGND VPWR VPWR __dut__.__uuf__._2215_/HI tie[160] sky130_fd_sc_hd__conb_1
XFILLER_102_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2400_ rst VGND VGND VPWR VPWR __dut__._2400_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2146_ VGND VGND VPWR VPWR __dut__.__uuf__._2146_/HI tie[91] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2077_ VGND VGND VPWR VPWR __dut__.__uuf__._2077_/HI tie[22] sky130_fd_sc_hd__conb_1
X__dut__._2331_ __dut__._2335_/A __dut__._2331_/B VGND VGND VPWR VPWR __dut__._2331_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2396__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2262_ __dut__._2262_/A1 __dut__._2262_/A2 __dut__._2261_/X VGND VGND VPWR
+ VPWR __dut__._2262_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1028_ __dut__.__uuf__._1241_/A __dut__._2227_/B __dut__._2225_/B
+ __dut__._2223_/B VGND VGND VPWR VPWR __dut__.__uuf__._1029_/D sky130_fd_sc_hd__or4_4
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2193_ __dut__._2213_/A __dut__._2193_/B VGND VGND VPWR VPWR __dut__._2193_/X
+ sky130_fd_sc_hd__and2_4
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_205 _242_/X VGND VGND VPWR VPWR psn_inst_psn_buff_339/A sky130_fd_sc_hd__buf_8
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_216 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1741_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_227 psn_inst_psn_buff_228/A VGND VGND VPWR VPWR __dut__._2355_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_129_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_249 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1729_/A
+ sky130_fd_sc_hd__buf_2
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_238 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2263_/A
+ sky130_fd_sc_hd__buf_2
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1977_ __dut__._2213_/A __dut__._1977_/B VGND VGND VPWR VPWR __dut__._1977_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_153_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1475__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2529_ rst VGND VGND VPWR VPWR __dut__._2529_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1488__A2 mp[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2000_ __dut__._1356_/X VGND VGND VPWR VPWR __dut__.__uuf__._2004_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_58_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1412__A2 mp[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1715_ __dut__._1959_/B __dut__._1969_/B VGND VGND VPWR VPWR __dut__.__uuf__._1716_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_147_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1646_ __dut__.__uuf__._1648_/A VGND VGND VPWR VPWR __dut__.__uuf__._1646_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2880_ __dut__._2892_/CLK __dut__._2880_/D __dut__._2372_/Y VGND VGND VPWR
+ VPWR __dut__._2880_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1900_ __dut__._1900_/A1 prod[7] __dut__._1899_/X VGND VGND VPWR VPWR __dut__._2869_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1831_ __dut__._1853_/A __dut__._2834_/Q VGND VGND VPWR VPWR __dut__._1831_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_135_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1577_ __dut__.__uuf__._1577_/A VGND VGND VPWR VPWR __dut__.__uuf__._1577_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1762_ __dut__._1854_/A1 tie[108] __dut__._1761_/X VGND VGND VPWR VPWR __dut__._2800_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1295__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1693_ __dut__._1693_/A __dut__._2765_/Q VGND VGND VPWR VPWR __dut__._1693_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2129_ VGND VGND VPWR VPWR __dut__.__uuf__._2129_/HI tie[74] sky130_fd_sc_hd__conb_1
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2314_ __dut__._2322_/A1 __dut__._2314_/A2 __dut__._2313_/X VGND VGND VPWR
+ VPWR __dut__._2314_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._1655__A __dut__.__uuf__._1655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_60_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2245_ __dut__._2251_/A __dut__._2245_/B VGND VGND VPWR VPWR __dut__._2245_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2176_ __dut__._2176_/A1 __dut__._2176_/A2 __dut__._2175_/X VGND VGND VPWR
+ VPWR __dut__._2176_/X sky130_fd_sc_hd__a21o_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1933__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1890__A2 prod[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_122_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2806__CLK clkbuf_opt_1_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1500_ __dut__.__uuf__._1516_/A VGND VGND VPWR VPWR __dut__.__uuf__._1500_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_144_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1431_ __dut__.__uuf__._1476_/A VGND VGND VPWR VPWR __dut__.__uuf__._1449_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_132_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1362_ __dut__.__uuf__._1711_/A VGND VGND VPWR VPWR __dut__.__uuf__._1362_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1293_ __dut__.__uuf__._1292_/Y __dut__.__uuf__._2047_/A __dut__.__uuf__._1283_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1293_/X sky130_fd_sc_hd__o21a_4
XFILLER_131_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1843__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2030_ __dut__._2030_/A1 __dut__._2030_/A2 __dut__._2029_/X VGND VGND VPWR
+ VPWR __dut__._2030_/X sky130_fd_sc_hd__a21o_4
XFILLER_26_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1629_ __dut__.__uuf__._1630_/A VGND VGND VPWR VPWR __dut__.__uuf__._1629_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2863_ _308_/CLK __dut__._2863_/D __dut__._2389_/Y VGND VGND VPWR VPWR __dut__._2863_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_135_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2794_ _270_/CLK __dut__._2794_/D __dut__._2458_/Y VGND VGND VPWR VPWR __dut__._2794_/Q
+ sky130_fd_sc_hd__dfrtp_4
X__dut__._1814_ __dut__._1854_/A1 tie[134] __dut__._1813_/X VGND VGND VPWR VPWR __dut__._2826_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_150_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1745_ __dut__._1745_/A __dut__._2791_/Q VGND VGND VPWR VPWR __dut__._1745_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_89_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1753__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1676_ __dut__._1726_/A1 tie[65] __dut__._1675_/X VGND VGND VPWR VPWR __dut__._2757_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_67_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2241__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2228_ __dut__._2228_/A1 __dut__._2228_/A2 __dut__._2227_/X VGND VGND VPWR
+ VPWR __dut__._2228_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2829__CLK __dut__._2845_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2584__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2159_ __dut__._2167_/A __dut__._2159_/B VGND VGND VPWR VPWR __dut__._2159_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1388__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1312__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_337_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1980_ __dut__._2059_/B __dut__._2065_/B __dut__.__uuf__._1979_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1981_/C sky130_fd_sc_hd__o21ai_4
XFILLER_63_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2494__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2394_ __dut__.__uuf__._2426_/CLK __dut__._2292_/X __dut__.__uuf__._1138_/X
+ VGND VGND VPWR VPWR __dut__._2293_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1414_ __dut__.__uuf__._1414_/A VGND VGND VPWR VPWR __dut__.__uuf__._1414_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1345_ __dut__.__uuf__._1342_/X __dut__.__uuf__._1344_/X __dut__._2191_/B
+ __dut__.__uuf__._1342_/X VGND VGND VPWR VPWR __dut__._2190_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1530_ __dut__._1530_/A1 __dut__._1528_/X __dut__._1529_/X VGND VGND VPWR
+ VPWR __dut__._2688_/D sky130_fd_sc_hd__a21o_4
XFILLER_113_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1573__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1276_ __dut__.__uuf__._1983_/A VGND VGND VPWR VPWR __dut__.__uuf__._1276_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1461_ __dut__._1461_/A __dut__._2660_/Q VGND VGND VPWR VPWR __dut__._1461_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_46_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1392_ __dut__._1282_/Y mp[2] __dut__._1391_/X VGND VGND VPWR VPWR __dut__._1392_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2013_ __dut__._2213_/A __dut__._2013_/B VGND VGND VPWR VPWR __dut__._2013_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_1 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1780_/A1 sky130_fd_sc_hd__buf_2
X_271_ _271_/CLK _271_/D VGND VGND VPWR VPWR _271_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_23_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2846_ clkbuf_opt_0_tck/X __dut__._2846_/D __dut__._2406_/Y VGND VGND VPWR
+ VPWR __dut__._2846_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2777_ __dut__._2869_/CLK __dut__._2777_/D __dut__._2475_/Y VGND VGND VPWR
+ VPWR __dut__._2777_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2579__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1728_ __dut__._1910_/A1 tie[91] __dut__._1727_/X VGND VGND VPWR VPWR __dut__._2783_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1483__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1659_ __dut__._1661_/A __dut__._2748_/Q VGND VGND VPWR VPWR __dut__._1659_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2651__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_287_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1130_ __dut__.__uuf__._1188_/A VGND VGND VPWR VPWR __dut__.__uuf__._1130_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2489__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2287__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_110_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1061_ __dut__.__uuf__._1071_/A VGND VGND VPWR VPWR __dut__.__uuf__._1061_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1963_ __dut__.__uuf__._1985_/A __dut__.__uuf__._1963_/B __dut__.__uuf__._1963_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1964_/A sky130_fd_sc_hd__or3_4
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1894_ __dut__.__uuf__._1894_/A VGND VGND VPWR VPWR __dut__.__uuf__._1894_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1772__A1 __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_30 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2014_/A1 sky130_fd_sc_hd__buf_2
XFILLER_152_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2700_ clkbuf_5_2_0_tck/X __dut__._2700_/D __dut__._2552_/Y VGND VGND VPWR
+ VPWR __dut__._2700_/Q sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_74 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2150_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_41 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2044_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_52 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2086_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_63 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2210_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_96 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1406_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._2631_ __dut__._2357_/B __dut__._2631_/D __dut__._2621_/Y VGND VGND VPWR
+ VPWR __dut__._2631_/Q sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_85 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1466_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1524__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2377_ __dut__.__uuf__._2412_/CLK __dut__._2258_/X __dut__.__uuf__._1187_/X
+ VGND VGND VPWR VPWR __dut__._2259_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2399__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2562_ rst VGND VGND VPWR VPWR __dut__._2562_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1328_ __dut__.__uuf__._1355_/A VGND VGND VPWR VPWR __dut__.__uuf__._1350_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2493_ rst VGND VGND VPWR VPWR __dut__._2493_/Y sky130_fd_sc_hd__inv_2
X__dut__._1513_ __dut__._1513_/A __dut__._2683_/Q VGND VGND VPWR VPWR __dut__._1513_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1259_ __dut__.__uuf__._1259_/A VGND VGND VPWR VPWR __dut__.__uuf__._1259_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1444_ __dut__._1282_/Y mp[14] __dut__._1443_/X VGND VGND VPWR VPWR __dut__._1444_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_86_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1375_ _234_/Y __dut__._2650_/Q VGND VGND VPWR VPWR __dut__._1375_/X sky130_fd_sc_hd__and2_4
XFILLER_27_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_254_ _308_/CLK _254_/D VGND VGND VPWR VPWR _255_/D sky130_fd_sc_hd__dfxtp_4
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_185_ _265_/Q _186_/B VGND VGND VPWR VPWR _264_/D sky130_fd_sc_hd__or2_4
XFILLER_142_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2829_ __dut__._2845_/CLK __dut__._2829_/D __dut__._2423_/Y VGND VGND VPWR
+ VPWR __dut__._2829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1941__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1754__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2300_ __dut__.__uuf__._2319_/CLK __dut__._2104_/X __dut__.__uuf__._1542_/X
+ VGND VGND VPWR VPWR __dut__._2105_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2231_ __dut__.__uuf__._2288_/CLK __dut__._1966_/X __dut__.__uuf__._1654_/X
+ VGND VGND VPWR VPWR __dut__._1967_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_125_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2162_ VGND VGND VPWR VPWR __dut__.__uuf__._2162_/HI tie[107] sky130_fd_sc_hd__conb_1
XFILLER_88_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2093_ VGND VGND VPWR VPWR __dut__.__uuf__._2093_/HI tie[38] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1113_ __dut__.__uuf__._1116_/A VGND VGND VPWR VPWR __dut__.__uuf__._1113_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1044_ __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR __dut__.__uuf__._2054_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1851__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1946_ __dut__._1336_/X VGND VGND VPWR VPWR __dut__.__uuf__._1950_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2302__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__306__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1877_ __dut__.__uuf__._1877_/A __dut__.__uuf__._1877_/B __dut__.__uuf__._1877_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1878_/A sky130_fd_sc_hd__or3_4
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1993_ __dut__._2213_/A __dut__._1993_/B VGND VGND VPWR VPWR __dut__._1993_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_124_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2614_ rst VGND VGND VPWR VPWR __dut__._2614_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2545_ rst VGND VGND VPWR VPWR __dut__._2545_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_90_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1580__A2 __dut__.__uuf__._1890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1761__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2476_ rst VGND VGND VPWR VPWR __dut__._2476_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1427_ _234_/Y __dut__._2663_/Q VGND VGND VPWR VPWR __dut__._1427_/X sky130_fd_sc_hd__and2_4
XFILLER_131_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1358_ __dut__._1358_/A1 __dut__._1356_/X __dut__._1357_/X VGND VGND VPWR
+ VPWR __dut__._2645_/D sky130_fd_sc_hd__a21o_4
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1289_ __dut__._1289_/A __dut__._2692_/Q VGND VGND VPWR VPWR __dut__._1289_/X
+ sky130_fd_sc_hd__and2_4
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_306_ _312_/CLK _306_/D trst VGND VGND VPWR VPWR _306_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2592__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_237_ _237_/A _297_/Q _300_/Q _237_/D VGND VGND VPWR VPWR _249_/D sky130_fd_sc_hd__or4_4
XFILLER_143_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_168_ _279_/Q _172_/B VGND VGND VPWR VPWR _278_/D sky130_fd_sc_hd__and2_4
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_152_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2325__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_65_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1800_ __dut__.__uuf__._1766_/X __dut__.__uuf__._1798_/B __dut__.__uuf__._1798_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1801_/C sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1731_ __dut__._1967_/B __dut__._1973_/B __dut__.__uuf__._1730_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1732_/C sky130_fd_sc_hd__o21ai_4
X__dut__.__uuf__._1662_ __dut__.__uuf__._2051_/A __dut__._1957_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1663_/A sky130_fd_sc_hd__and2_4
XFILLER_119_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2007__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1593_ __dut__.__uuf__._1593_/A VGND VGND VPWR VPWR __dut__.__uuf__._1593_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_106_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2214_ VGND VGND VPWR VPWR __dut__.__uuf__._2214_/HI tie[159] sky130_fd_sc_hd__conb_1
XANTENNA___dut__.__uuf__._1478__A __dut__.__uuf__._1478_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2145_ VGND VGND VPWR VPWR __dut__.__uuf__._2145_/HI tie[90] sky130_fd_sc_hd__conb_1
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2076_ VGND VGND VPWR VPWR __dut__.__uuf__._2076_/HI tie[21] sky130_fd_sc_hd__conb_1
X__dut__._2330_ __dut__._2338_/A1 __dut__._2330_/A2 __dut__._2329_/X VGND VGND VPWR
+ VPWR __dut__._2330_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2261_ __dut__._2261_/A __dut__._2261_/B VGND VGND VPWR VPWR __dut__._2261_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1027_ __dut__._2229_/B VGND VGND VPWR VPWR __dut__.__uuf__._1241_/A
+ sky130_fd_sc_hd__inv_2
X__dut__._2192_ __dut__._2200_/A1 __dut__._2192_/A2 __dut__._2191_/X VGND VGND VPWR
+ VPWR __dut__._2192_/X sky130_fd_sc_hd__a21o_4
XFILLER_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_206 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR psn_inst_psn_buff_208/A
+ sky130_fd_sc_hd__buf_2
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_217 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2337_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_228 psn_inst_psn_buff_228/A VGND VGND VPWR VPWR __dut__._2349_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_101_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_239 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2261_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1929_ __dut__.__uuf__._1983_/A VGND VGND VPWR VPWR __dut__.__uuf__._1929_/X
+ sky130_fd_sc_hd__buf_2
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2862__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1718__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1976_ __dut__._2078_/A1 __dut__._1976_/A2 __dut__._1975_/X VGND VGND VPWR
+ VPWR __dut__._1976_/X sky130_fd_sc_hd__a21o_4
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1388__A __dut__.__uuf__._1711_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2587__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2528_ rst VGND VGND VPWR VPWR __dut__._2528_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__299__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1491__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2459_ rst VGND VGND VPWR VPWR __dut__._2459_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1298__A __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2497__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1714_ __dut__._1284_/X VGND VGND VPWR VPWR __dut__.__uuf__._1718_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_119_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1645_ __dut__.__uuf__._1648_/A VGND VGND VPWR VPWR __dut__.__uuf__._1645_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1830_ __dut__._1854_/A1 tie[142] __dut__._1829_/X VGND VGND VPWR VPWR __dut__._2834_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1576_ __dut__.__uuf__._1564_/X __dut__.__uuf__._1559_/X __dut__._2089_/B
+ __dut__.__uuf__._1462_/A __dut__.__uuf__._1575_/X VGND VGND VPWR VPWR __dut__._2088_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_135_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1761_ __dut__._1853_/A __dut__._2799_/Q VGND VGND VPWR VPWR __dut__._1761_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_103_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1692_ __dut__._1694_/A1 tie[73] __dut__._1691_/X VGND VGND VPWR VPWR __dut__._2765_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2128_ VGND VGND VPWR VPWR __dut__.__uuf__._2128_/HI tie[73] sky130_fd_sc_hd__conb_1
XFILLER_57_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2059_ VGND VGND VPWR VPWR __dut__.__uuf__._2059_/HI tie[4] sky130_fd_sc_hd__conb_1
X__dut__._2313_ __dut__._2313_/A __dut__._2313_/B VGND VGND VPWR VPWR __dut__._2313_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2244_ __dut__._2244_/A1 __dut__._2244_/A2 __dut__._2243_/X VGND VGND VPWR
+ VPWR __dut__._2244_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2175_ __dut__._2189_/A __dut__._2175_/B VGND VGND VPWR VPWR __dut__._2175_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_53_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1959_ __dut__._2213_/A __dut__._1959_/B VGND VGND VPWR VPWR __dut__._1959_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_97_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_115_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1430_ __dut__.__uuf__._1418_/X __dut__.__uuf__._1428_/X __dut__._2157_/B
+ __dut__.__uuf__._1429_/X VGND VGND VPWR VPWR __dut__._2156_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1361_ __dut__._2185_/B VGND VGND VPWR VPWR __dut__.__uuf__._1361_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_132_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1292_ __dut__._2211_/B VGND VGND VPWR VPWR __dut__.__uuf__._1292_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_86_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_tck clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR clkbuf_3_7_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_54_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1628_ __dut__.__uuf__._1630_/A VGND VGND VPWR VPWR __dut__.__uuf__._1628_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2346__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2862_ _308_/CLK __dut__._2862_/D __dut__._2390_/Y VGND VGND VPWR VPWR __dut__._2862_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_135_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2793_ _270_/CLK __dut__._2793_/D __dut__._2459_/Y VGND VGND VPWR VPWR __dut__._2793_/Q
+ sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1559_ __dut__.__uuf__._1578_/A VGND VGND VPWR VPWR __dut__.__uuf__._1559_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1813_ __dut__._1813_/A __dut__._2825_/Q VGND VGND VPWR VPWR __dut__._1813_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1744_ __dut__._1854_/A1 tie[99] __dut__._1743_/X VGND VGND VPWR VPWR __dut__._2791_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_150_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1675_ __dut__._1701_/A __dut__._2756_/Q VGND VGND VPWR VPWR __dut__._1675_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_83_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2227_ __dut__._2227_/A __dut__._2227_/B VGND VGND VPWR VPWR __dut__._2227_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_83_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0___dut__.__uuf__.__clk_source__ clkbuf_4_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2282_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__._2158_ __dut__._2166_/A1 __dut__._2158_/A2 __dut__._2157_/X VGND VGND VPWR
+ VPWR __dut__._2158_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1388__A2 mp[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2089_ __dut__._2095_/A __dut__._2089_/B VGND VGND VPWR VPWR __dut__._2089_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_145_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1312__A2 mc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_232_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1413_ __dut__.__uuf__._1711_/A VGND VGND VPWR VPWR __dut__.__uuf__._1413_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_144_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2393_ __dut__.__uuf__._2415_/CLK __dut__._2290_/X __dut__.__uuf__._1140_/X
+ VGND VGND VPWR VPWR __dut__._2291_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_117_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1344_ __dut__.__uuf__._1343_/Y __dut__.__uuf__._1336_/X __dut__.__uuf__._1337_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1344_/X sky130_fd_sc_hd__o21a_4
XFILLER_132_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1275_ __dut__.__uuf__._1765_/A VGND VGND VPWR VPWR __dut__.__uuf__._1983_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_100_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1460_ __dut__._1282_/Y mc[4] __dut__._1459_/X VGND VGND VPWR VPWR __dut__._1460_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1391_ _234_/Y __dut__._2654_/Q VGND VGND VPWR VPWR __dut__._1391_/X sky130_fd_sc_hd__and2_4
XFILLER_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2012_ __dut__._2012_/A1 __dut__._2012_/A2 __dut__._2011_/X VGND VGND VPWR
+ VPWR __dut__._2012_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_2 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1778_/A1 sky130_fd_sc_hd__buf_2
XFILLER_139_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_270_ _270_/CLK _270_/D VGND VGND VPWR VPWR _270_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_16_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2845_ __dut__._2845_/CLK __dut__._2845_/D __dut__._2407_/Y VGND VGND VPWR
+ VPWR __dut__._2845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2776_ __dut__._2869_/CLK __dut__._2776_/D __dut__._2476_/Y VGND VGND VPWR
+ VPWR __dut__._2776_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1727_ __dut__._1729_/A __dut__._2782_/Q VGND VGND VPWR VPWR __dut__._1727_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1658_ __dut__._1658_/A1 tie[56] __dut__._1657_/X VGND VGND VPWR VPWR __dut__._2748_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1589_ __dut__._1793_/A __dut__._2713_/Q VGND VGND VPWR VPWR __dut__._1589_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2595__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1939__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_182_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1060_ __dut__.__uuf__._2054_/A VGND VGND VPWR VPWR __dut__.__uuf__._1071_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_95_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1962_ __dut__.__uuf__._1929_/X __dut__.__uuf__._1960_/B __dut__.__uuf__._1960_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1963_/C sky130_fd_sc_hd__o21a_4
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1893_ __dut__._2027_/B __dut__._2033_/B VGND VGND VPWR VPWR __dut__.__uuf__._1894_/A
+ sky130_fd_sc_hd__and2_4
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1849__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_20 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1860_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_31 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2024_/A1 sky130_fd_sc_hd__buf_2
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_42 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1330_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_64 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2214_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_53 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2084_/A1 sky130_fd_sc_hd__buf_2
XFILLER_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2376_ __dut__.__uuf__._2412_/CLK __dut__._2256_/X __dut__.__uuf__._1190_/X
+ VGND VGND VPWR VPWR __dut__._2257_/B sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_86 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1450_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_97 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1402_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._2630_ __dut__._2357_/B __dut__._2630_/D __dut__._2622_/Y VGND VGND VPWR
+ VPWR __dut__._2630_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1524__A2 start VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_75 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2228_/A1 sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1327_ __dut__.__uuf__._1315_/X __dut__.__uuf__._1325_/X __dut__._2197_/B
+ __dut__.__uuf__._1326_/X VGND VGND VPWR VPWR __dut__._2196_/A2 sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__.__uuf__._2231__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_132_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2561_ rst VGND VGND VPWR VPWR __dut__._2561_/Y sky130_fd_sc_hd__inv_2
X__dut__._2492_ rst VGND VGND VPWR VPWR __dut__._2492_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1288__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1512_ __dut__._1282_/Y mp[29] __dut__._1511_/X VGND VGND VPWR VPWR __dut__._1512_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1258_ __dut__.__uuf__._1269_/A VGND VGND VPWR VPWR __dut__.__uuf__._1258_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1443_ _234_/Y __dut__._2667_/Q VGND VGND VPWR VPWR __dut__._1443_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1189_ __dut__.__uuf__._1177_/X __dut__.__uuf__._1188_/X __dut__._2259_/B
+ __dut__._2261_/B __dut__.__uuf__._1185_/X VGND VGND VPWR VPWR __dut__._2258_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_73_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1944__A __dut__.__uuf__._1998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1374_ __dut__._2044_/A1 __dut__._1372_/X __dut__._1373_/X VGND VGND VPWR
+ VPWR __dut__._2649_/D sky130_fd_sc_hd__a21o_4
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1460__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1759__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_253_ _308_/CLK tms VGND VGND VPWR VPWR _254_/D sky130_fd_sc_hd__dfxtp_4
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_184_ _266_/Q _186_/B VGND VGND VPWR VPWR _265_/D sky130_fd_sc_hd__or2_4
XFILLER_127_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2828_ _193_/A __dut__._2828_/D __dut__._2424_/Y VGND VGND VPWR VPWR __dut__._2828_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_151_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2759_ __dut__._2767_/CLK __dut__._2759_/D __dut__._2493_/Y VGND VGND VPWR
+ VPWR __dut__._2759_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2230_ __dut__.__uuf__._2355_/CLK __dut__._1964_/X __dut__.__uuf__._1656_/X
+ VGND VGND VPWR VPWR __dut__._1965_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_130_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2161_ VGND VGND VPWR VPWR __dut__.__uuf__._2161_/HI tie[106] sky130_fd_sc_hd__conb_1
XFILLER_88_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2092_ VGND VGND VPWR VPWR __dut__.__uuf__._2092_/HI tie[37] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1112_ __dut__.__uuf__._1103_/X __dut__.__uuf__._1100_/X __dut__._2311_/B
+ __dut__._2313_/B __dut__.__uuf__._1111_/X VGND VGND VPWR VPWR __dut__._2310_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1043_ __dut__.__uuf__._1089_/A VGND VGND VPWR VPWR __dut__.__uuf__._1618_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_110_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1945_ __dut__.__uuf__._1937_/A __dut__.__uuf__._1942_/B __dut__.__uuf__._1944_/X
+ VGND VGND VPWR VPWR __dut__._2042_/A2 sky130_fd_sc_hd__o21a_4
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1876_ __dut__.__uuf__._1875_/X __dut__.__uuf__._1873_/B __dut__.__uuf__._1873_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1877_/C sky130_fd_sc_hd__o21a_4
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1579__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1992_ __dut__._2000_/A1 __dut__._1992_/A2 __dut__._1991_/X VGND VGND VPWR
+ VPWR __dut__._1992_/X sky130_fd_sc_hd__a21o_4
XFILLER_124_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2613_ rst VGND VGND VPWR VPWR __dut__._2613_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2359_ __dut__.__uuf__._2402_/CLK __dut__._2222_/X __dut__.__uuf__._1258_/X
+ VGND VGND VPWR VPWR __dut__._2223_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2203__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2544_ rst VGND VGND VPWR VPWR __dut__._2544_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_83_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2475_ rst VGND VGND VPWR VPWR __dut__._2475_/Y sky130_fd_sc_hd__inv_2
X__dut__._1426_ __dut__._1426_/A1 __dut__._1424_/X __dut__._1425_/X VGND VGND VPWR
+ VPWR __dut__._2662_/D sky130_fd_sc_hd__a21o_4
XFILLER_62_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1357_ __dut__._1361_/A __dut__._2644_/Q VGND VGND VPWR VPWR __dut__._1357_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1288_ __dut__._1282_/Y mc[10] __dut__._1287_/X VGND VGND VPWR VPWR __dut__._1288_/X
+ sky130_fd_sc_hd__a21o_4
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_305_ _312_/CLK _305_/D trst VGND VGND VPWR VPWR _305_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_236_ _236_/A _236_/B _298_/Q _236_/D VGND VGND VPWR VPWR _237_/D sky130_fd_sc_hd__and4_4
X_167_ _280_/Q _172_/B VGND VGND VPWR VPWR _279_/D sky130_fd_sc_hd__and2_4
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2113__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_145_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_312_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1424__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1730_ __dut__.__uuf__._1730_/A VGND VGND VPWR VPWR __dut__.__uuf__._1730_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1399__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1661_ __dut__.__uuf__._2054_/A VGND VGND VPWR VPWR __dut__.__uuf__._1661_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1592_ __dut__.__uuf__._1593_/A VGND VGND VPWR VPWR __dut__.__uuf__._1592_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2213_ VGND VGND VPWR VPWR __dut__.__uuf__._2213_/HI tie[158] sky130_fd_sc_hd__conb_1
XFILLER_115_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2144_ VGND VGND VPWR VPWR __dut__.__uuf__._2144_/HI tie[89] sky130_fd_sc_hd__conb_1
XFILLER_130_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2075_ VGND VGND VPWR VPWR __dut__.__uuf__._2075_/HI tie[20] sky130_fd_sc_hd__conb_1
Xclkbuf_5_9_0_tck clkbuf_5_9_0_tck/A VGND VGND VPWR VPWR clkbuf_5_9_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2260_ __dut__._2260_/A1 __dut__._2260_/A2 __dut__._2259_/X VGND VGND VPWR
+ VPWR __dut__._2260_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1026_ __dut__._2219_/B VGND VGND VPWR VPWR __dut__.__uuf__._1234_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_71_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2191_ __dut__._2213_/A __dut__._2191_/B VGND VGND VPWR VPWR __dut__._2191_/X
+ sky130_fd_sc_hd__and2_4
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_207 psn_inst_psn_buff_208/A VGND VGND VPWR VPWR __dut__._1745_/A
+ sky130_fd_sc_hd__buf_2
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_218 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2335_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1928_ __dut__.__uuf__._1928_/A VGND VGND VPWR VPWR __dut__.__uuf__._1931_/B
+ sky130_fd_sc_hd__inv_2
Xpsn_inst_psn_buff_229 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2269_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_101_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1859_ __dut__._1300_/X VGND VGND VPWR VPWR __dut__.__uuf__._1863_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_138_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1975_ __dut__._2213_/A __dut__._1975_/B VGND VGND VPWR VPWR __dut__._1975_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_153_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2527_ rst VGND VGND VPWR VPWR __dut__._2527_/Y sky130_fd_sc_hd__inv_2
X__dut__._2458_ rst VGND VGND VPWR VPWR __dut__._2458_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1409_ __dut__._1433_/A __dut__._2657_/Q VGND VGND VPWR VPWR __dut__._1409_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2389_ rst VGND VGND VPWR VPWR __dut__._2389_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_219_ _219_/A _224_/B VGND VGND VPWR VPWR _292_/D sky130_fd_sc_hd__and2_4
XFILLER_128_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1947__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_262_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1948__A2 prod[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1713_ __dut__.__uuf__._1966_/A VGND VGND VPWR VPWR __dut__.__uuf__._1742_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_119_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1644_ __dut__.__uuf__._1648_/A VGND VGND VPWR VPWR __dut__.__uuf__._1644_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1857__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1575_ __dut__._1388_/X __dut__.__uuf__._1565_/X __dut__._2091_/B
+ __dut__.__uuf__._1309_/A VGND VGND VPWR VPWR __dut__.__uuf__._1575_/X sky130_fd_sc_hd__o22a_4
XFILLER_135_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1760_ __dut__._1854_/A1 tie[107] __dut__._1759_/X VGND VGND VPWR VPWR __dut__._2799_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_150_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1691_ __dut__._1691_/A __dut__._2764_/Q VGND VGND VPWR VPWR __dut__._1691_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_102_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2127_ VGND VGND VPWR VPWR __dut__.__uuf__._2127_/HI tie[72] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2058_ VGND VGND VPWR VPWR __dut__.__uuf__._2058_/HI tie[3] sky130_fd_sc_hd__conb_1
X__dut__._2312_ __dut__._2322_/A1 __dut__._2312_/A2 __dut__._2311_/X VGND VGND VPWR
+ VPWR __dut__._2312_/X sky130_fd_sc_hd__a21o_4
XANTENNA__253__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_tck tck VGND VGND VPWR VPWR clkbuf_0_tck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_44_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2243_ __dut__._2243_/A __dut__._2243_/B VGND VGND VPWR VPWR __dut__._2243_/X
+ sky130_fd_sc_hd__and2_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2174_ __dut__._2176_/A1 __dut__._2174_/A2 __dut__._2173_/X VGND VGND VPWR
+ VPWR __dut__._2174_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_46_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1767__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2315__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_137_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1958_ __dut__._1958_/A1 __dut__._1958_/A2 __dut__._1957_/X VGND VGND VPWR
+ VPWR __dut__._1958_/X sky130_fd_sc_hd__a21o_4
XFILLER_140_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1889_ __dut__._2313_/A __dut__._2863_/Q VGND VGND VPWR VPWR __dut__._1889_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2598__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_108_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1360_ __dut__.__uuf__._1375_/A VGND VGND VPWR VPWR __dut__.__uuf__._1360_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1291_ __dut__.__uuf__._1295_/A VGND VGND VPWR VPWR __dut__.__uuf__._1291_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2852__CLK clkbuf_5_6_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2301__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2861_ _193_/A __dut__._2861_/D __dut__._2391_/Y VGND VGND VPWR VPWR _209_/A2
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1587__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1627_ __dut__.__uuf__._1630_/A VGND VGND VPWR VPWR __dut__.__uuf__._1627_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1812_ __dut__._1854_/A1 tie[133] __dut__._1811_/X VGND VGND VPWR VPWR __dut__._2825_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2792_ _193_/A __dut__._2792_/D __dut__._2460_/Y VGND VGND VPWR VPWR __dut__._2792_/Q
+ sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1558_ __dut__.__uuf__._1558_/A VGND VGND VPWR VPWR __dut__.__uuf__._1558_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_122_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1743_ __dut__._1743_/A __dut__._2790_/Q VGND VGND VPWR VPWR __dut__._1743_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1489_ __dut__._1480_/X __dut__.__uuf__._1480_/X __dut__._2133_/B
+ __dut__.__uuf__._1485_/X VGND VGND VPWR VPWR __dut__.__uuf__._1489_/X sky130_fd_sc_hd__o22a_4
XFILLER_107_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1674_ __dut__._1726_/A1 tie[64] __dut__._1673_/X VGND VGND VPWR VPWR __dut__._2756_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_131_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._2211__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2282__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2226_ __dut__._2228_/A1 __dut__._2226_/A2 __dut__._2225_/X VGND VGND VPWR
+ VPWR __dut__._2226_/X sky130_fd_sc_hd__a21o_4
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2157_ __dut__._2167_/A __dut__._2157_/B VGND VGND VPWR VPWR __dut__._2157_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2088_ __dut__._2088_/A1 __dut__._2088_/A2 __dut__._2087_/X VGND VGND VPWR
+ VPWR __dut__._2088_/X sky130_fd_sc_hd__a21o_4
XFILLER_9_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1848__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2121__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1784__B1 __dut__._1783_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1412_ __dut__._2165_/B VGND VGND VPWR VPWR __dut__.__uuf__._1412_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2392_ __dut__.__uuf__._2426_/CLK __dut__._2288_/X __dut__.__uuf__._1143_/X
+ VGND VGND VPWR VPWR __dut__._2289_/B sky130_fd_sc_hd__dfrtp_4
Xclkbuf_4_15_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2422_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_144_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1343_ __dut__._2193_/B VGND VGND VPWR VPWR __dut__.__uuf__._1343_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_144_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1274_ __dut__._2215_/B VGND VGND VPWR VPWR __dut__.__uuf__._1765_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_113_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1390_ __dut__._1390_/A1 __dut__._1388_/X __dut__._1389_/X VGND VGND VPWR
+ VPWR __dut__._2653_/D sky130_fd_sc_hd__a21o_4
XFILLER_39_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2011_ __dut__._2213_/A __dut__._2011_/B VGND VGND VPWR VPWR __dut__._2011_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_42_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_3 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1776_/A1 sky130_fd_sc_hd__buf_2
XFILLER_139_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2844_ __dut__._2845_/CLK __dut__._2844_/D __dut__._2408_/Y VGND VGND VPWR
+ VPWR __dut__._2844_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2775_ __dut__._2869_/CLK __dut__._2775_/D __dut__._2477_/Y VGND VGND VPWR
+ VPWR __dut__._2775_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1726_ __dut__._1726_/A1 tie[90] __dut__._1725_/X VGND VGND VPWR VPWR __dut__._2782_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_77_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1657_ __dut__._1661_/A __dut__._2747_/Q VGND VGND VPWR VPWR __dut__._1657_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1588_ __dut__._1790_/A1 tie[21] __dut__._1587_/X VGND VGND VPWR VPWR __dut__._2713_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_91_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2209_ __dut__._2213_/A __dut__._2209_/B VGND VGND VPWR VPWR __dut__._2209_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1766__B1 __dut__._1765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_tck clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR clkbuf_3_5_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_142_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1587__A __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_175_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1961_ __dut__.__uuf__._1961_/A VGND VGND VPWR VPWR __dut__.__uuf__._1963_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1892_ __dut__._1312_/X VGND VGND VPWR VPWR __dut__.__uuf__._1896_/B
+ sky130_fd_sc_hd__inv_2
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_10 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1880_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_21 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1858_/A1 sky130_fd_sc_hd__buf_2
XFILLER_117_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_43 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1378_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_32 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2016_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_65 __dut__._1772_/A1 VGND VGND VPWR VPWR psn_inst_psn_buff_73/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_54 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2080_/A1 sky130_fd_sc_hd__buf_2
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1865__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_87 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2112_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_98 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1398_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2375_ __dut__.__uuf__._2412_/CLK __dut__._2254_/X __dut__.__uuf__._1195_/X
+ VGND VGND VPWR VPWR __dut__._2255_/B sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_76 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2146_/A1 sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1041__B1 __dut__._1961_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1326_ __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR __dut__.__uuf__._1326_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_99_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2560_ rst VGND VGND VPWR VPWR __dut__._2560_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1288__A2 mc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2491_ rst VGND VGND VPWR VPWR __dut__._2491_/Y sky130_fd_sc_hd__inv_2
X__dut__._1511_ _234_/Y __dut__._2684_/Q VGND VGND VPWR VPWR __dut__._1511_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1257_ __dut__.__uuf__._1255_/Y __dut__.__uuf__._1256_/X __dut__.__uuf__._1229_/X
+ __dut__._2225_/B __dut__.__uuf__._1247_/X VGND VGND VPWR VPWR __dut__._2224_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_104_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1442_ __dut__._1442_/A1 __dut__._1440_/X __dut__._1441_/X VGND VGND VPWR
+ VPWR __dut__._2666_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1188_ __dut__.__uuf__._1188_/A VGND VGND VPWR VPWR __dut__.__uuf__._1188_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1373_ __dut__._2095_/A __dut__._2638_/Q VGND VGND VPWR VPWR __dut__._1373_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2846__D __dut__._2846_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1460__A2 mc[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_252_ _198_/A _305_/Q VGND VGND VPWR VPWR _252_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ _267_/Q _190_/B VGND VGND VPWR VPWR _266_/D sky130_fd_sc_hd__and2_4
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1775__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2827_ _308_/CLK __dut__._2827_/D __dut__._2425_/Y VGND VGND VPWR VPWR __dut__._2827_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2758_ __dut__._2767_/CLK __dut__._2758_/D __dut__._2494_/Y VGND VGND VPWR
+ VPWR __dut__._2758_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1200__A __dut__.__uuf__._1215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1709_ __dut__._1709_/A __dut__._2773_/Q VGND VGND VPWR VPWR __dut__._1709_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2689_ clkbuf_5_3_0_tck/X __dut__._2689_/D __dut__._2563_/Y VGND VGND VPWR
+ VPWR __dut__._2689_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_292_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_1_0___dut__.__uuf__.__clk_source___A clkbuf_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2160_ VGND VGND VPWR VPWR __dut__.__uuf__._2160_/HI tie[105] sky130_fd_sc_hd__conb_1
XFILLER_141_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2091_ VGND VGND VPWR VPWR __dut__.__uuf__._2091_/HI tie[36] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1111_ __dut__.__uuf__._1141_/A VGND VGND VPWR VPWR __dut__.__uuf__._1111_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_96_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1042_ rst VGND VGND VPWR VPWR __dut__.__uuf__._1089_/A sky130_fd_sc_hd__inv_2
XFILLER_141_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1944_ __dut__.__uuf__._1998_/A VGND VGND VPWR VPWR __dut__.__uuf__._1944_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_51_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1875_ __dut__.__uuf__._1983_/A VGND VGND VPWR VPWR __dut__.__uuf__._1875_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_137_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1991_ __dut__._2213_/A __dut__._1991_/B VGND VGND VPWR VPWR __dut__._1991_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1595__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2612_ rst VGND VGND VPWR VPWR __dut__._2612_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2358_ __dut__.__uuf__._2398_/CLK __dut__._2220_/X __dut__.__uuf__._1262_/X
+ VGND VGND VPWR VPWR __dut__._2221_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_78_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2543_ rst VGND VGND VPWR VPWR __dut__._2543_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1309_ __dut__.__uuf__._1309_/A VGND VGND VPWR VPWR __dut__.__uuf__._1309_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2289_ __dut__.__uuf__._2355_/CLK __dut__._2082_/X __dut__.__uuf__._1583_/X
+ VGND VGND VPWR VPWR __dut__._2083_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2474_ rst VGND VGND VPWR VPWR __dut__._2474_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_76_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1425_ __dut__._1433_/A __dut__._2661_/Q VGND VGND VPWR VPWR __dut__._1425_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_131_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1356_ __dut__._1282_/Y mc[26] __dut__._1355_/X VGND VGND VPWR VPWR __dut__._1356_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1287_ _234_/Y __dut__._2628_/Q VGND VGND VPWR VPWR __dut__._1287_/X sky130_fd_sc_hd__and2_4
XFILLER_15_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_304_ _308_/CLK _304_/D trst VGND VGND VPWR VPWR _304_/Q sky130_fd_sc_hd__dfstp_4
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_235_ _235_/A _311_/Q VGND VGND VPWR VPWR _236_/D sky130_fd_sc_hd__nor2_4
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_166_ _281_/Q _171_/B VGND VGND VPWR VPWR _280_/D sky130_fd_sc_hd__or2_4
XFILLER_6_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_138_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1424__A2 mp[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2809__CLK clkbuf_opt_1_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_psn_inst_psn_buff_305_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1660_ __dut__.__uuf__._1660_/A VGND VGND VPWR VPWR __dut__.__uuf__._1660_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1591_ __dut__.__uuf__._1593_/A VGND VGND VPWR VPWR __dut__.__uuf__._1591_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_146_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2212_ VGND VGND VPWR VPWR __dut__.__uuf__._2212_/HI tie[157] sky130_fd_sc_hd__conb_1
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2143_ VGND VGND VPWR VPWR __dut__.__uuf__._2143_/HI tie[88] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._1360__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2074_ VGND VGND VPWR VPWR __dut__.__uuf__._2074_/HI tie[19] sky130_fd_sc_hd__conb_1
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1025_ __dut__._1955_/B VGND VGND VPWR VPWR __dut__.__uuf__._2051_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2190_ __dut__._2200_/A1 __dut__._2190_/A2 __dut__._2189_/X VGND VGND VPWR
+ VPWR __dut__._2190_/X sky130_fd_sc_hd__a21o_4
XFILLER_45_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_208 psn_inst_psn_buff_208/A VGND VGND VPWR VPWR __dut__._1853_/A
+ sky130_fd_sc_hd__buf_8
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_219 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2273_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1927_ __dut__.__uuf__._1960_/A __dut__.__uuf__._1927_/B __dut__.__uuf__._1927_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1928_/A sky130_fd_sc_hd__or3_4
XFILLER_101_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1858_ __dut__.__uuf__._1966_/A VGND VGND VPWR VPWR __dut__.__uuf__._1906_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1789_ __dut__.__uuf__._1789_/A VGND VGND VPWR VPWR __dut__.__uuf__._1791_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_125_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1974_ __dut__._2078_/A1 __dut__._1974_/A2 __dut__._1973_/X VGND VGND VPWR
+ VPWR __dut__._1974_/X sky130_fd_sc_hd__a21o_4
XFILLER_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2526_ rst VGND VGND VPWR VPWR __dut__._2526_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2457_ rst VGND VGND VPWR VPWR __dut__._2457_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2244__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1408_ __dut__._1282_/Y mp[6] __dut__._1407_/X VGND VGND VPWR VPWR __dut__._1408_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._2388_ rst VGND VGND VPWR VPWR __dut__._2388_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1339_ _234_/Y __dut__._2641_/Q VGND VGND VPWR VPWR __dut__._1339_/X sky130_fd_sc_hd__and2_4
XFILLER_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_218_ _292_/Q _291_/Q _217_/X VGND VGND VPWR VPWR _291_/D sky130_fd_sc_hd__o21a_4
XFILLER_144_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_149_ _145_/Y _294_/Q _306_/Q _305_/Q _219_/A VGND VGND VPWR VPWR _305_/D sky130_fd_sc_hd__o32a_4
XFILLER_143_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1963__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_255_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1712_ __dut__.__uuf__._1765_/A VGND VGND VPWR VPWR __dut__.__uuf__._1966_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1643_ __dut__.__uuf__._1643_/A VGND VGND VPWR VPWR __dut__.__uuf__._1648_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1574_ __dut__.__uuf__._1577_/A VGND VGND VPWR VPWR __dut__.__uuf__._1574_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1873__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1690_ __dut__._1690_/A1 tie[72] __dut__._1689_/X VGND VGND VPWR VPWR __dut__._2764_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2126_ VGND VGND VPWR VPWR __dut__.__uuf__._2126_/HI tie[71] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2057_ VGND VGND VPWR VPWR __dut__.__uuf__._2057_/HI tie[2] sky130_fd_sc_hd__conb_1
X__dut__._2311_ __dut__._2313_/A __dut__._2311_/B VGND VGND VPWR VPWR __dut__._2311_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_17_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2242_ __dut__._2244_/A1 __dut__._2242_/A2 __dut__._2241_/X VGND VGND VPWR
+ VPWR __dut__._2242_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2173_ __dut__._2189_/A __dut__._2173_/B VGND VGND VPWR VPWR __dut__._2173_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_44_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2209__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_39_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1957_ __dut__._2213_/A __dut__._1957_/B VGND VGND VPWR VPWR __dut__._1957_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_140_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1783__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1324__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1888_ __dut__._2356_/A1 prod[1] __dut__._1887_/X VGND VGND VPWR VPWR __dut__._2863_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_97_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2509_ rst VGND VGND VPWR VPWR __dut__._2509_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2119__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__304__SET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_8_0_tck clkbuf_5_9_0_tck/A VGND VGND VPWR VPWR clkbuf_5_8_0_tck/X sky130_fd_sc_hd__clkbuf_1
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1290_ __dut__.__uuf__._1286_/X __dut__.__uuf__._1289_/X __dut__._2211_/B
+ __dut__.__uuf__._1286_/X VGND VGND VPWR VPWR __dut__._2210_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2860_ clkbuf_5_5_0_tck/X __dut__._2860_/D __dut__._2392_/Y VGND VGND VPWR
+ VPWR __dut__._2860_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1626_ __dut__.__uuf__._1630_/A VGND VGND VPWR VPWR __dut__.__uuf__._1626_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1557_ __dut__.__uuf__._1543_/X __dut__.__uuf__._1538_/X __dut__._2099_/B
+ __dut__.__uuf__._1548_/X __dut__.__uuf__._1556_/X VGND VGND VPWR VPWR __dut__._2098_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1811_ __dut__._1811_/A __dut__._2824_/Q VGND VGND VPWR VPWR __dut__._1811_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_107_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2791_ _312_/CLK __dut__._2791_/D __dut__._2461_/Y VGND VGND VPWR VPWR __dut__._2791_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_122_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1488_ __dut__.__uuf__._1494_/A VGND VGND VPWR VPWR __dut__.__uuf__._1488_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1742_ __dut__._1854_/A1 tie[98] __dut__._1741_/X VGND VGND VPWR VPWR __dut__._2790_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1673_ __dut__._1673_/A __dut__._2755_/Q VGND VGND VPWR VPWR __dut__._1673_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_103_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2109_ VGND VGND VPWR VPWR __dut__.__uuf__._2109_/HI tie[54] sky130_fd_sc_hd__conb_1
XFILLER_123_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2225_ __dut__._2227_/A __dut__._2225_/B VGND VGND VPWR VPWR __dut__._2225_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2156_ __dut__._2166_/A1 __dut__._2156_/A2 __dut__._2155_/X VGND VGND VPWR
+ VPWR __dut__._2156_/X sky130_fd_sc_hd__a21o_4
X__dut__._2087_ __dut__._2213_/A __dut__._2087_/B VGND VGND VPWR VPWR __dut__._2087_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1203__A __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2402__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2034__A __dut__.__uuf__._2044_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_120_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_218_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1536__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1411_ __dut__.__uuf__._1426_/A VGND VGND VPWR VPWR __dut__.__uuf__._1411_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2391_ __dut__.__uuf__._2426_/CLK __dut__._2286_/X __dut__.__uuf__._1146_/X
+ VGND VGND VPWR VPWR __dut__._2287_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1342_ __dut__.__uuf__._1393_/A VGND VGND VPWR VPWR __dut__.__uuf__._1342_/X
+ sky130_fd_sc_hd__buf_2
Xclkbuf_3_7_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0___dut__.__uuf__.__clk_source__/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1273_ __dut__.__uuf__._1295_/A VGND VGND VPWR VPWR __dut__.__uuf__._1273_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2305__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2010_ __dut__._2010_/A1 __dut__._2010_/A2 __dut__._2009_/X VGND VGND VPWR
+ VPWR __dut__._2010_/X sky130_fd_sc_hd__a21o_4
XFILLER_42_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_4 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1774_/A1 sky130_fd_sc_hd__buf_2
XFILLER_139_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1609_ __dut__.__uuf__._1611_/A VGND VGND VPWR VPWR __dut__.__uuf__._1609_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2843_ clkbuf_opt_2_tck/A __dut__._2843_/D __dut__._2409_/Y VGND VGND VPWR
+ VPWR __dut__._2843_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2774_ __dut__._2869_/CLK __dut__._2774_/D __dut__._2478_/Y VGND VGND VPWR
+ VPWR __dut__._2774_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1725_ __dut__._1729_/A __dut__._2781_/Q VGND VGND VPWR VPWR __dut__._1725_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1656_ __dut__._1658_/A1 tie[55] __dut__._1655_/X VGND VGND VPWR VPWR __dut__._2747_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1587_ __dut__._1793_/A __dut__._2712_/Q VGND VGND VPWR VPWR __dut__._1587_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2208_ __dut__._2208_/A1 __dut__._2208_/A2 __dut__._2207_/X VGND VGND VPWR
+ VPWR __dut__._2208_/X sky130_fd_sc_hd__a21o_4
XANTENNA__266__CLK _270_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2139_ __dut__._2149_/A __dut__._2139_/B VGND VGND VPWR VPWR __dut__._2139_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_9_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2842__CLK clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1971__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_168_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_335_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1960_ __dut__.__uuf__._1960_/A __dut__.__uuf__._1960_/B __dut__.__uuf__._1960_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1961_/A sky130_fd_sc_hd__or3_4
XFILLER_36_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1891_ __dut__.__uuf__._1883_/A __dut__.__uuf__._1888_/B __dut__.__uuf__._1890_/X
+ VGND VGND VPWR VPWR __dut__._2022_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_149_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2307__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_11 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1878_/A1 sky130_fd_sc_hd__buf_2
XFILLER_136_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_22 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1856_/A1 sky130_fd_sc_hd__buf_2
XFILLER_117_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_44 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1286_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_33 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2008_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_55 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2082_/A1 sky130_fd_sc_hd__buf_2
XFILLER_155_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_88 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1446_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_99 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2110_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2374_ __dut__.__uuf__._2412_/CLK __dut__._2252_/X __dut__.__uuf__._1197_/X
+ VGND VGND VPWR VPWR __dut__._2253_/B sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_77 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2144_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_66 psn_inst_psn_buff_73/A VGND VGND VPWR VPWR __dut__._2152_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1041__B2 __dut__.__uuf__._1040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1325_ __dut__.__uuf__._1324_/Y __dut__.__uuf__._1309_/X __dut__.__uuf__._1311_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1325_/X sky130_fd_sc_hd__o21a_4
XFILLER_120_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1510_ __dut__._1510_/A1 __dut__._1508_/X __dut__._1509_/X VGND VGND VPWR
+ VPWR __dut__._2683_/D sky130_fd_sc_hd__a21o_4
X__dut__._2490_ rst VGND VGND VPWR VPWR __dut__._2490_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1256_ __dut__._2225_/B __dut__.__uuf__._1259_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1256_/X sky130_fd_sc_hd__or2_4
XANTENNA___dut__._1881__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1187_ __dut__.__uuf__._1190_/A VGND VGND VPWR VPWR __dut__.__uuf__._1187_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1441_ __dut__._1441_/A __dut__._2665_/Q VGND VGND VPWR VPWR __dut__._1441_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1372_ __dut__._1282_/Y mc[2] __dut__._1371_/X VGND VGND VPWR VPWR __dut__._1372_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__243__A1 tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1748__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_251_ _195_/X _257_/Q VGND VGND VPWR VPWR _251_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_psn_inst_psn_buff_21_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_182_ _182_/A VGND VGND VPWR VPWR _190_/B sky130_fd_sc_hd__buf_2
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2826_ _308_/CLK __dut__._2826_/D __dut__._2426_/Y VGND VGND VPWR VPWR __dut__._2826_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_123_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2757_ __dut__._2767_/CLK __dut__._2757_/D __dut__._2495_/Y VGND VGND VPWR
+ VPWR __dut__._2757_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1708_ __dut__._1726_/A1 tie[81] __dut__._1707_/X VGND VGND VPWR VPWR __dut__._2773_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2688_ __dut__._2894_/CLK __dut__._2688_/D __dut__._2564_/Y VGND VGND VPWR
+ VPWR __dut__._2688_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1639_ __dut__._1661_/A __dut__._2738_/Q VGND VGND VPWR VPWR __dut__._1639_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1791__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2127__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_285_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1110_ __dut__.__uuf__._1116_/A VGND VGND VPWR VPWR __dut__.__uuf__._1110_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2090_ VGND VGND VPWR VPWR __dut__.__uuf__._2090_/HI tie[35] sky130_fd_sc_hd__conb_1
XFILLER_56_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1041_ __dut__.__uuf__._1034_/X __dut__.__uuf__._1038_/X __dut__._1885_/B
+ __dut__._1961_/B __dut__.__uuf__._1040_/X VGND VGND VPWR VPWR __dut__._2356_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1943_ __dut__.__uuf__._1943_/A VGND VGND VPWR VPWR __dut__._2044_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_34_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1874_ __dut__.__uuf__._1874_/A VGND VGND VPWR VPWR __dut__.__uuf__._1877_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_149_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1990_ __dut__._2000_/A1 __dut__._1990_/A2 __dut__._1989_/X VGND VGND VPWR
+ VPWR __dut__._1990_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2426_ __dut__.__uuf__._2426_/CLK __dut__._2356_/X __dut__.__uuf__._2054_/X
+ VGND VGND VPWR VPWR __dut__._1885_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_79_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2611_ rst VGND VGND VPWR VPWR __dut__._2611_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2357_ __dut__.__uuf__._2398_/CLK __dut__._2218_/X __dut__.__uuf__._1265_/X
+ VGND VGND VPWR VPWR __dut__._2219_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_120_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2542_ rst VGND VGND VPWR VPWR __dut__._2542_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1308_ __dut__.__uuf__._1771_/A VGND VGND VPWR VPWR __dut__.__uuf__._1309_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2288_ __dut__.__uuf__._2288_/CLK __dut__._2080_/X __dut__.__uuf__._1584_/X
+ VGND VGND VPWR VPWR __dut__._2081_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2500__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1239_ __dut__._2227_/B __dut__.__uuf__._1255_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1242_/B sky130_fd_sc_hd__and2_4
XFILLER_115_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2473_ rst VGND VGND VPWR VPWR __dut__._2473_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1424_ __dut__._1282_/Y mp[9] __dut__._1423_/X VGND VGND VPWR VPWR __dut__._1424_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1355_ _234_/Y __dut__._2645_/Q VGND VGND VPWR VPWR __dut__._1355_/X sky130_fd_sc_hd__and2_4
Xclkbuf_2_1_0_tck clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR clkbuf_3_3_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_131_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1286_ __dut__._1286_/A1 __dut__._1284_/X __dut__._1285_/X VGND VGND VPWR
+ VPWR __dut__._2627_/D sky130_fd_sc_hd__a21o_4
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_303_ _303_/CLK _303_/D trst VGND VGND VPWR VPWR _303_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_234_ _304_/Q VGND VGND VPWR VPWR _234_/Y sky130_fd_sc_hd__inv_4
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_165_ _282_/Q _172_/B VGND VGND VPWR VPWR _281_/D sky130_fd_sc_hd__and2_4
XFILLER_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__304__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2809_ clkbuf_opt_1_tck/X __dut__._2809_/D __dut__._2443_/Y VGND VGND VPWR
+ VPWR __dut__._2809_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2410__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1590_ __dut__.__uuf__._1593_/A VGND VGND VPWR VPWR __dut__.__uuf__._1590_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2211_ VGND VGND VPWR VPWR __dut__.__uuf__._2211_/HI tie[156] sky130_fd_sc_hd__conb_1
XFILLER_142_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2142_ VGND VGND VPWR VPWR __dut__.__uuf__._2142_/HI tie[87] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._1360__A2 mc[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2073_ VGND VGND VPWR VPWR __dut__.__uuf__._2073_/HI tie[18] sky130_fd_sc_hd__conb_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_209 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1743_/A
+ sky130_fd_sc_hd__buf_2
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1820__B1 __dut__._1819_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1926_ __dut__._2039_/B __dut__._2045_/B __dut__.__uuf__._1925_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1927_/C sky130_fd_sc_hd__o21ai_4
XFILLER_61_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1857_ __dut__.__uuf__._1850_/A __dut__.__uuf__._1855_/B __dut__.__uuf__._1836_/X
+ VGND VGND VPWR VPWR __dut__._2010_/A2 sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1788_ __dut__.__uuf__._1798_/A __dut__.__uuf__._1788_/B __dut__.__uuf__._1788_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1789_/A sky130_fd_sc_hd__or3_4
XFILLER_137_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1973_ __dut__._2213_/A __dut__._1973_/B VGND VGND VPWR VPWR __dut__._1973_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_133_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2409_ __dut__.__uuf__._2412_/CLK __dut__._2322_/X __dut__.__uuf__._1094_/X
+ VGND VGND VPWR VPWR __dut__._2323_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_121_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2525_ rst VGND VGND VPWR VPWR __dut__._2525_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2456_ rst VGND VGND VPWR VPWR __dut__._2456_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2300__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1407_ _234_/Y __dut__._2658_/Q VGND VGND VPWR VPWR __dut__._1407_/X sky130_fd_sc_hd__and2_4
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2387_ rst VGND VGND VPWR VPWR __dut__._2387_/Y sky130_fd_sc_hd__inv_2
X__dut__._1338_ __dut__._1346_/A1 __dut__._1336_/X __dut__._1337_/X VGND VGND VPWR
+ VPWR __dut__._2640_/D sky130_fd_sc_hd__a21o_4
XFILLER_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_217_ _229_/A VGND VGND VPWR VPWR _217_/X sky130_fd_sc_hd__buf_2
XFILLER_11_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2405__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_148_ _237_/A _141_/Y _307_/Q _306_/Q _143_/Y VGND VGND VPWR VPWR _306_/D sky130_fd_sc_hd__a32o_4
XFILLER_98_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_opt_2_tck_A clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_150_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_248_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0___dut__.__uuf__.__clk_source__ clkbuf_2_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1711_ __dut__.__uuf__._1711_/A VGND VGND VPWR VPWR __dut__.__uuf__._1768_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1642_ __dut__.__uuf__._1642_/A VGND VGND VPWR VPWR __dut__.__uuf__._1642_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2358__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1573_ __dut__.__uuf__._1564_/X __dut__.__uuf__._1559_/X __dut__._2091_/B
+ __dut__.__uuf__._1462_/A __dut__.__uuf__._1572_/X VGND VGND VPWR VPWR __dut__._2090_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_147_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2125_ VGND VGND VPWR VPWR __dut__.__uuf__._2125_/HI tie[70] sky130_fd_sc_hd__conb_1
XFILLER_102_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2056_ VGND VGND VPWR VPWR __dut__.__uuf__._2056_/HI tie[1] sky130_fd_sc_hd__conb_1
X__dut__._2310_ __dut__._2356_/A1 __dut__._2310_/A2 __dut__._2309_/X VGND VGND VPWR
+ VPWR __dut__._2310_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2241_ __dut__._2243_/A __dut__._2241_/B VGND VGND VPWR VPWR __dut__._2241_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_112_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2172_ __dut__._2176_/A1 __dut__._2172_/A2 __dut__._2171_/X VGND VGND VPWR
+ VPWR __dut__._2172_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1909_ __dut__.__uuf__._1931_/A __dut__.__uuf__._1909_/B __dut__.__uuf__._1909_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1910_/A sky130_fd_sc_hd__or3_4
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1956_ __dut__._2228_/A1 __dut__._1956_/A2 __dut__._1955_/X VGND VGND VPWR
+ VPWR __dut__._1956_/X sky130_fd_sc_hd__a21o_4
XFILLER_141_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1783__B __dut__._2810_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1324__A2 mc[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1887_ __dut__._2313_/A __dut__._2862_/Q VGND VGND VPWR VPWR __dut__._1887_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1696__A __dut__._1528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2508_ rst VGND VGND VPWR VPWR __dut__._2508_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2361__CLK __dut__.__uuf__._2402_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_62_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2439_ rst VGND VGND VPWR VPWR __dut__._2439_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2135__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1625_ __dut__.__uuf__._1643_/A VGND VGND VPWR VPWR __dut__.__uuf__._1630_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_135_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1810_ __dut__._1810_/A1 tie[132] __dut__._1809_/X VGND VGND VPWR VPWR __dut__._2824_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1556_ __dut__._1408_/X __dut__.__uuf__._1544_/X __dut__._2101_/B
+ __dut__.__uuf__._1549_/X VGND VGND VPWR VPWR __dut__.__uuf__._1556_/X sky130_fd_sc_hd__o22a_4
XFILLER_123_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2234__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2790_ _312_/CLK __dut__._2790_/D __dut__._2462_/Y VGND VGND VPWR VPWR __dut__._2790_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_89_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1487_ __dut__.__uuf__._1478_/X __dut__.__uuf__._1473_/X __dut__._2133_/B
+ __dut__.__uuf__._1484_/X __dut__.__uuf__._1486_/X VGND VGND VPWR VPWR __dut__._2132_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1741_ __dut__._1741_/A __dut__._2789_/Q VGND VGND VPWR VPWR __dut__._1741_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1672_ __dut__._1672_/A1 tie[63] __dut__._1671_/X VGND VGND VPWR VPWR __dut__._2755_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__310__SET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2108_ VGND VGND VPWR VPWR __dut__.__uuf__._2108_/HI tie[53] sky130_fd_sc_hd__conb_1
XFILLER_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2039_ __dut__.__uuf__._2032_/A __dut__.__uuf__._2037_/B __dut__.__uuf__._1998_/X
+ VGND VGND VPWR VPWR __dut__._2078_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_123_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2224_ __dut__._2228_/A1 __dut__._2224_/A2 __dut__._2223_/X VGND VGND VPWR
+ VPWR __dut__._2224_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_51_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2155_ __dut__._2167_/A __dut__._2155_/B VGND VGND VPWR VPWR __dut__._2155_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2086_ __dut__._2086_/A1 __dut__._2086_/A2 __dut__._2085_/X VGND VGND VPWR
+ VPWR __dut__._2086_/X sky130_fd_sc_hd__a21o_4
XFILLER_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1939_ __dut__._2327_/A __dut__._2888_/Q VGND VGND VPWR VPWR __dut__._1939_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1969__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_113_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__292__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1536__A2 mc[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2390_ __dut__.__uuf__._2426_/CLK __dut__._2284_/X __dut__.__uuf__._1150_/X
+ VGND VGND VPWR VPWR __dut__._2285_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1410_ __dut__.__uuf__._1404_/X __dut__.__uuf__._1409_/X __dut__._2165_/B
+ __dut__.__uuf__._1404_/X VGND VGND VPWR VPWR __dut__._2164_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1341_ __dut__.__uuf__._1341_/A VGND VGND VPWR VPWR __dut__.__uuf__._1393_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_144_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1272_ __dut__.__uuf__._1355_/A VGND VGND VPWR VPWR __dut__.__uuf__._1295_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1472__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1879__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpsn_inst_psn_buff_5 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1770_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__309__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1608_ __dut__.__uuf__._1611_/A VGND VGND VPWR VPWR __dut__.__uuf__._1608_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2842_ clkbuf_opt_2_tck/A __dut__._2842_/D __dut__._2410_/Y VGND VGND VPWR
+ VPWR __dut__._2842_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2773_ __dut__._2869_/CLK __dut__._2773_/D __dut__._2479_/Y VGND VGND VPWR
+ VPWR __dut__._2773_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2503__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1539_ __dut__._1428_/X __dut__.__uuf__._1523_/X __dut__._2109_/B
+ __dut__.__uuf__._1528_/X VGND VGND VPWR VPWR __dut__.__uuf__._1539_/X sky130_fd_sc_hd__o22a_4
XFILLER_150_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2794__CLK _270_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1724_ __dut__._1726_/A1 tie[89] __dut__._1723_/X VGND VGND VPWR VPWR __dut__._2781_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_89_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_99_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1655_ __dut__._1661_/A __dut__._2746_/Q VGND VGND VPWR VPWR __dut__._1655_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1586_ __dut__._1790_/A1 tie[20] __dut__._1585_/X VGND VGND VPWR VPWR __dut__._2712_/D
+ sky130_fd_sc_hd__a21o_4
Xclkbuf_5_7_0_tck clkbuf_5_7_0_tck/A VGND VGND VPWR VPWR clkbuf_opt_1_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_94_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2207_ __dut__._2213_/A __dut__._2207_/B VGND VGND VPWR VPWR __dut__._2207_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1789__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2138_ __dut__._2140_/A1 __dut__._2138_/A2 __dut__._2137_/X VGND VGND VPWR
+ VPWR __dut__._2138_/X sky130_fd_sc_hd__a21o_4
X__dut__._2069_ __dut__._2213_/A __dut__._2069_/B VGND VGND VPWR VPWR __dut__._2069_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2413__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_230_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_328_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1890_ __dut__.__uuf__._1890_/A VGND VGND VPWR VPWR __dut__.__uuf__._1890_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_118_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_12 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1876_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_23 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1806_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_34 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2010_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_45 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1382_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_56 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1958_/A1 sky130_fd_sc_hd__buf_2
XFILLER_145_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_89 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1442_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2373_ __dut__.__uuf__._2412_/CLK __dut__._2250_/X __dut__.__uuf__._1199_/X
+ VGND VGND VPWR VPWR __dut__._2251_/B sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_78 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2136_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_67 psn_inst_psn_buff_73/A VGND VGND VPWR VPWR __dut__._2154_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1041__A2 __dut__.__uuf__._1038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1324_ __dut__._2199_/B VGND VGND VPWR VPWR __dut__.__uuf__._1324_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1255_ __dut__.__uuf__._1255_/A VGND VGND VPWR VPWR __dut__.__uuf__._1255_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_101_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1440_ __dut__._1282_/Y mp[13] __dut__._1439_/X VGND VGND VPWR VPWR __dut__._1440_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1186_ __dut__.__uuf__._1177_/X __dut__.__uuf__._1174_/X __dut__._2261_/B
+ __dut__._2263_/B __dut__.__uuf__._1185_/X VGND VGND VPWR VPWR __dut__._2260_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_104_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1371_ _234_/Y __dut__._2649_/Q VGND VGND VPWR VPWR __dut__._1371_/X sky130_fd_sc_hd__and2_4
XFILLER_39_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_250_ _196_/X _313_/Q VGND VGND VPWR VPWR _250_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_181_ _268_/Q _181_/B VGND VGND VPWR VPWR _267_/D sky130_fd_sc_hd__and2_4
XFILLER_129_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_14_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2233__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2825_ _308_/CLK __dut__._2825_/D __dut__._2427_/Y VGND VGND VPWR VPWR __dut__._2825_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2756_ __dut__._2767_/CLK __dut__._2756_/D __dut__._2496_/Y VGND VGND VPWR
+ VPWR __dut__._2756_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1707_ __dut__._1707_/A __dut__._2772_/Q VGND VGND VPWR VPWR __dut__._1707_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2687_ __dut__._2894_/CLK __dut__._2687_/D __dut__._2565_/Y VGND VGND VPWR
+ VPWR __dut__._2687_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1638_ __dut__._1658_/A1 tie[46] __dut__._1637_/X VGND VGND VPWR VPWR __dut__._2738_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1569_ __dut__._1611_/A __dut__._2703_/Q VGND VGND VPWR VPWR __dut__._1569_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1209__A __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1436__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2408__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0___dut__.__uuf__.__clk_source__ clkbuf_4_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2278_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__.__uuf__._1271__A2 __dut__.__uuf__._1040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._2143__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_180_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_278_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1040_ __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR __dut__.__uuf__._1040_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_83_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1942_ __dut__.__uuf__._1985_/A __dut__.__uuf__._1942_/B __dut__.__uuf__._1942_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1943_/A sky130_fd_sc_hd__or3_4
XFILLER_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1873_ __dut__.__uuf__._1906_/A __dut__.__uuf__._1873_/B __dut__.__uuf__._1873_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1874_/A sky130_fd_sc_hd__or3_4
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._2053__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2425_ __dut__.__uuf__._2426_/CLK __dut__._2354_/X __dut__.__uuf__._1057_/A
+ VGND VGND VPWR VPWR __dut__._2355_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_117_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2610_ rst VGND VGND VPWR VPWR __dut__._2610_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1902__A2 prod[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2356_ __dut__.__uuf__._2398_/CLK __dut__._2216_/X __dut__.__uuf__._1269_/X
+ VGND VGND VPWR VPWR __dut__._2217_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_105_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2541_ rst VGND VGND VPWR VPWR __dut__._2541_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1307_ __dut__.__uuf__._1307_/A VGND VGND VPWR VPWR __dut__.__uuf__._1771_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2287_ __dut__.__uuf__._2323_/CLK __dut__._2078_/X __dut__.__uuf__._1585_/X
+ VGND VGND VPWR VPWR __dut__._2079_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_120_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2472_ rst VGND VGND VPWR VPWR __dut__._2472_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1238_ __dut__._2225_/B __dut__.__uuf__._1259_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1255_/A sky130_fd_sc_hd__and2_4
XANTENNA__256__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1423_ _234_/Y __dut__._2662_/Q VGND VGND VPWR VPWR __dut__._1423_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2832__CLK __dut__._2845_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1169_ __dut__.__uuf__._1162_/X __dut__.__uuf__._1159_/X __dut__._2273_/B
+ __dut__._2275_/B __dut__.__uuf__._1156_/X VGND VGND VPWR VPWR __dut__._2272_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1354_ __dut__._1354_/A1 __dut__._1352_/X __dut__._1353_/X VGND VGND VPWR
+ VPWR __dut__._2644_/D sky130_fd_sc_hd__a21o_4
XFILLER_55_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1285_ tdi __dut__._2313_/A VGND VGND VPWR VPWR __dut__._1285_/X sky130_fd_sc_hd__and2_4
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ _303_/CLK _302_/D trst VGND VGND VPWR VPWR _302_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_233_ _249_/Q VGND VGND VPWR VPWR tdo_paden_o sky130_fd_sc_hd__inv_2
XFILLER_156_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2318__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_164_ _182_/A VGND VGND VPWR VPWR _172_/B sky130_fd_sc_hd__buf_2
XFILLER_7_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2808_ clkbuf_opt_1_tck/A __dut__._2808_/D __dut__._2444_/Y VGND VGND VPWR
+ VPWR __dut__._2808_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2739_ __dut__._2894_/CLK __dut__._2739_/D __dut__._2513_/Y VGND VGND VPWR
+ VPWR __dut__._2739_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1307__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1977__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2210_ VGND VGND VPWR VPWR __dut__.__uuf__._2210_/HI tie[155] sky130_fd_sc_hd__conb_1
XFILLER_114_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2855__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2141_ VGND VGND VPWR VPWR __dut__.__uuf__._2141_/HI tie[86] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2601__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2072_ VGND VGND VPWR VPWR __dut__.__uuf__._2072_/HI tie[17] sky130_fd_sc_hd__conb_1
XFILLER_68_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1925_ __dut__.__uuf__._1925_/A VGND VGND VPWR VPWR __dut__.__uuf__._1925_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1820__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1856_ __dut__.__uuf__._1856_/A VGND VGND VPWR VPWR __dut__._2012_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1787_ __dut__._1987_/B __dut__._1993_/B __dut__.__uuf__._1786_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1788_/C sky130_fd_sc_hd__o21ai_4
XANTENNA___dut__._1887__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1972_ __dut__._2078_/A1 __dut__._1972_/A2 __dut__._1971_/X VGND VGND VPWR
+ VPWR __dut__._1972_/X sky130_fd_sc_hd__a21o_4
XFILLER_152_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2408_ __dut__.__uuf__._2412_/CLK __dut__._2320_/X __dut__.__uuf__._1096_/X
+ VGND VGND VPWR VPWR __dut__._2321_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1031__B __dut__._1957_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2511__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2339_ __dut__.__uuf__._2348_/CLK __dut__._2182_/X __dut__.__uuf__._1360_/X
+ VGND VGND VPWR VPWR __dut__._2183_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_121_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2524_ rst VGND VGND VPWR VPWR __dut__._2524_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_81_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2455_ rst VGND VGND VPWR VPWR __dut__._2455_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1406_ __dut__._1406_/A1 __dut__._1404_/X __dut__._1405_/X VGND VGND VPWR
+ VPWR __dut__._2657_/D sky130_fd_sc_hd__a21o_4
X__dut__._2386_ rst VGND VGND VPWR VPWR __dut__._2386_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1337_ __dut__._1341_/A __dut__._2639_/Q VGND VGND VPWR VPWR __dut__._1337_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_31_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1797__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_216_ _291_/Q _231_/A VGND VGND VPWR VPWR _290_/D sky130_fd_sc_hd__and2_4
X_147_ _307_/Q _145_/Y _294_/Q _146_/X VGND VGND VPWR VPWR _307_/D sky130_fd_sc_hd__a211o_4
XANTENNA___dut__.__uuf__._2290__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_144_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2421__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_143_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_310_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1710_ __dut__._1885_/B __dut__.__uuf__._1681_/A __dut__._2293_/B
+ __dut__.__uuf__._1682_/A VGND VGND VPWR VPWR prod[31] sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1641_ __dut__.__uuf__._1642_/A VGND VGND VPWR VPWR __dut__.__uuf__._1641_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2358__A2 clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1572_ __dut__._1392_/X __dut__.__uuf__._1565_/X __dut__._2093_/B
+ __dut__.__uuf__._1309_/A VGND VGND VPWR VPWR __dut__.__uuf__._1572_/X sky130_fd_sc_hd__o22a_4
XFILLER_134_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_tck clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR clkbuf_3_1_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_143_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2124_ VGND VGND VPWR VPWR __dut__.__uuf__._2124_/HI tie[69] sky130_fd_sc_hd__conb_1
XFILLER_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2055_ VGND VGND VPWR VPWR __dut__.__uuf__._2055_/HI tie[0] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2294__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2240_ __dut__._2244_/A1 __dut__._2240_/A2 __dut__._2239_/X VGND VGND VPWR
+ VPWR __dut__._2240_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2171_ __dut__._2189_/A __dut__._2171_/B VGND VGND VPWR VPWR __dut__._2171_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1908_ __dut__.__uuf__._1875_/X __dut__.__uuf__._1906_/B __dut__.__uuf__._1906_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1909_/C sky130_fd_sc_hd__o21a_4
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1839_ __dut__._2007_/B __dut__._2013_/B VGND VGND VPWR VPWR __dut__.__uuf__._1840_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_40_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2506__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__.__uuf__._1042__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1955_ __dut__._2147_/A __dut__._1955_/B VGND VGND VPWR VPWR __dut__._1955_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_137_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1886_ __dut__._2356_/A1 prod[0] __dut__._1885_/X VGND VGND VPWR VPWR __dut__._2862_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2507_ rst VGND VGND VPWR VPWR __dut__._2507_/Y sky130_fd_sc_hd__inv_2
X__dut__._2438_ rst VGND VGND VPWR VPWR __dut__._2438_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2369_ rst VGND VGND VPWR VPWR __dut__._2369_/Y sky130_fd_sc_hd__inv_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2416__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2151__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_260_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1624_ __dut__.__uuf__._1624_/A VGND VGND VPWR VPWR __dut__.__uuf__._1624_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1555_ __dut__.__uuf__._1558_/A VGND VGND VPWR VPWR __dut__.__uuf__._1555_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1740_ __dut__._2328_/A1 tie[97] __dut__._1739_/X VGND VGND VPWR VPWR __dut__._2789_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1486_ __dut__._1484_/X __dut__.__uuf__._1480_/X __dut__._2135_/B
+ __dut__.__uuf__._1485_/X VGND VGND VPWR VPWR __dut__.__uuf__._1486_/X sky130_fd_sc_hd__o22a_4
XFILLER_131_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1671_ __dut__._1673_/A __dut__._2754_/Q VGND VGND VPWR VPWR __dut__._1671_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2061__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2107_ VGND VGND VPWR VPWR __dut__.__uuf__._2107_/HI tie[52] sky130_fd_sc_hd__conb_1
Xclkbuf_opt_0_tck clkbuf_opt_1_tck/A VGND VGND VPWR VPWR clkbuf_opt_0_tck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2038_ __dut__.__uuf__._2038_/A VGND VGND VPWR VPWR __dut__._2080_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2223_ __dut__._2227_/A __dut__._2223_/B VGND VGND VPWR VPWR __dut__._2223_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_60_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__.__uuf__._1037__A __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2154_ __dut__._2154_/A1 __dut__._2154_/A2 __dut__._2153_/X VGND VGND VPWR
+ VPWR __dut__._2154_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_44_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_opt_1_tck_A clkbuf_opt_1_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2085_ __dut__._2213_/A __dut__._2085_/B VGND VGND VPWR VPWR __dut__._2085_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_154_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1938_ __dut__._2328_/A1 prod[26] __dut__._1937_/X VGND VGND VPWR VPWR __dut__._2888_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1869_ __dut__._2213_/A __dut__._2853_/Q VGND VGND VPWR VPWR __dut__._1869_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_107_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1315__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_106_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1985__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1340_ __dut__.__uuf__._1350_/A VGND VGND VPWR VPWR __dut__.__uuf__._1340_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_113_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1271_ __dut__._2217_/B __dut__.__uuf__._1040_/X __dut__.__uuf__._1234_/B
+ __dut__.__uuf__._1270_/X VGND VGND VPWR VPWR __dut__._2216_/A2 sky130_fd_sc_hd__o22a_4
XFILLER_112_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1472__A2 mp[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_6 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1768_/A1 sky130_fd_sc_hd__buf_2
XFILLER_147_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1607_ __dut__.__uuf__._1611_/A VGND VGND VPWR VPWR __dut__.__uuf__._1607_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2841_ clkbuf_opt_2_tck/A __dut__._2841_/D __dut__._2411_/Y VGND VGND VPWR
+ VPWR __dut__._2841_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__.__uuf__._2351__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2772_ __dut__._2869_/CLK __dut__._2772_/D __dut__._2480_/Y VGND VGND VPWR
+ VPWR __dut__._2772_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1538_ __dut__.__uuf__._1578_/A VGND VGND VPWR VPWR __dut__.__uuf__._1538_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1723_ __dut__._1729_/A __dut__._2780_/Q VGND VGND VPWR VPWR __dut__._1723_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1469_ __dut__.__uuf__._1472_/A VGND VGND VPWR VPWR __dut__.__uuf__._1469_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1654_ __dut__._1658_/A1 tie[54] __dut__._1653_/X VGND VGND VPWR VPWR __dut__._2746_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_77_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1585_ __dut__._1793_/A __dut__._2711_/Q VGND VGND VPWR VPWR __dut__._1585_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2206_ __dut__._2206_/A1 __dut__._2206_/A2 __dut__._2205_/X VGND VGND VPWR
+ VPWR __dut__._2206_/X sky130_fd_sc_hd__a21o_4
X__dut__._2137_ __dut__._2149_/A __dut__._2137_/B VGND VGND VPWR VPWR __dut__._2137_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2068_ __dut__._2068_/A1 __dut__._2068_/A2 __dut__._2067_/X VGND VGND VPWR
+ VPWR __dut__._2068_/X sky130_fd_sc_hd__a21o_4
XFILLER_139_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_190 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2248_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_13 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1874_/A1 sky130_fd_sc_hd__buf_2
XFILLER_118_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_24 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1804_/A1 sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2604__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_46 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1386_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_35 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2012_/A1 sky130_fd_sc_hd__buf_2
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2372_ __dut__.__uuf__._2372_/CLK __dut__._2248_/X __dut__.__uuf__._1202_/X
+ VGND VGND VPWR VPWR __dut__._2249_/B sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_79 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2140_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_57 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1964_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_68 psn_inst_psn_buff_73/A VGND VGND VPWR VPWR __dut__._2184_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1323_ __dut__.__uuf__._1323_/A VGND VGND VPWR VPWR __dut__.__uuf__._1323_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1254_ __dut__.__uuf__._1269_/A VGND VGND VPWR VPWR __dut__.__uuf__._1254_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1185_ __dut__.__uuf__._1215_/A VGND VGND VPWR VPWR __dut__.__uuf__._1185_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1370_ __dut__._1378_/A1 __dut__._1368_/X __dut__._1369_/X VGND VGND VPWR
+ VPWR __dut__._2648_/D sky130_fd_sc_hd__a21o_4
XFILLER_104_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1315__A __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_180_ _269_/Q _181_/B VGND VGND VPWR VPWR _268_/D sky130_fd_sc_hd__and2_4
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2514__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2824_ clkbuf_5_1_0_tck/X __dut__._2824_/D __dut__._2428_/Y VGND VGND VPWR
+ VPWR __dut__._2824_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__.__uuf__._1050__A __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2755_ __dut__._2767_/CLK __dut__._2755_/D __dut__._2497_/Y VGND VGND VPWR
+ VPWR __dut__._2755_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1706_ __dut__._1726_/A1 tie[80] __dut__._1705_/X VGND VGND VPWR VPWR __dut__._2772_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2686_ __dut__._2744_/CLK __dut__._2686_/D __dut__._2566_/Y VGND VGND VPWR
+ VPWR __dut__._2686_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1637_ __dut__._1661_/A __dut__._2737_/Q VGND VGND VPWR VPWR __dut__._1637_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1568_ __dut__._1568_/A1 tie[11] __dut__._1567_/X VGND VGND VPWR VPWR __dut__._2703_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2247__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_92_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1499_ _234_/Y __dut__._2681_/Q VGND VGND VPWR VPWR __dut__._1499_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1436__A2 mp[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2424__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1372__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_173_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1941_ __dut__.__uuf__._1929_/X __dut__.__uuf__._1939_/B __dut__.__uuf__._1939_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1942_/C sky130_fd_sc_hd__o21a_4
XFILLER_24_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1503__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1872_ __dut__._2019_/B __dut__._2025_/B __dut__.__uuf__._1871_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1873_/C sky130_fd_sc_hd__o21ai_4
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_6_0_tck clkbuf_5_7_0_tck/A VGND VGND VPWR VPWR clkbuf_5_6_0_tck/X sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2424_ __dut__.__uuf__._2426_/CLK __dut__._2352_/X __dut__.__uuf__._1047_/X
+ VGND VGND VPWR VPWR __dut__._2353_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_11_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2415_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2355_ __dut__.__uuf__._2355_/CLK __dut__._2214_/X __dut__.__uuf__._1273_/X
+ VGND VGND VPWR VPWR __dut__._2215_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1306_ __dut__._2205_/B VGND VGND VPWR VPWR __dut__.__uuf__._1306_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_132_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2540_ rst VGND VGND VPWR VPWR __dut__._2540_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2286_ __dut__.__uuf__._2288_/CLK __dut__._2076_/X __dut__.__uuf__._1586_/X
+ VGND VGND VPWR VPWR __dut__._2077_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2471_ rst VGND VGND VPWR VPWR __dut__._2471_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1237_ __dut__._2223_/B __dut__.__uuf__._1260_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1259_/A sky130_fd_sc_hd__and2_4
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1422_ __dut__._1422_/A1 __dut__._1420_/X __dut__._1421_/X VGND VGND VPWR
+ VPWR __dut__._2661_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1168_ __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR __dut__.__uuf__._1168_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1353_ __dut__._1361_/A __dut__._2643_/Q VGND VGND VPWR VPWR __dut__._1353_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1099_ __dut__.__uuf__._1102_/A VGND VGND VPWR VPWR __dut__.__uuf__._1099_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_39_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2509__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1284_ mc[0] __dut__._1282_/Y __dut__._1283_/X VGND VGND VPWR VPWR __dut__._1284_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_301_ _312_/CLK _301_/D trst VGND VGND VPWR VPWR _301_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1045__A __dut__.__uuf__._2054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_232_ _304_/Q _231_/B _217_/X VGND VGND VPWR VPWR _303_/D sky130_fd_sc_hd__o21a_4
XFILLER_156_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_163_ _283_/Q _163_/B VGND VGND VPWR VPWR _282_/D sky130_fd_sc_hd__and2_4
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2807_ clkbuf_opt_1_tck/A __dut__._2807_/D __dut__._2445_/Y VGND VGND VPWR
+ VPWR __dut__._2807_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2738_ __dut__._2744_/CLK __dut__._2738_/D __dut__._2514_/Y VGND VGND VPWR
+ VPWR __dut__._2738_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2669_ __dut__._2680_/CLK __dut__._2669_/D __dut__._2583_/Y VGND VGND VPWR
+ VPWR __dut__._2669_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2419__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1323__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_290_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1993__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1896__A2 prod[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2140_ VGND VGND VPWR VPWR __dut__.__uuf__._2140_/HI tie[85] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2071_ VGND VGND VPWR VPWR __dut__.__uuf__._2071_/HI tie[16] sky130_fd_sc_hd__conb_1
XFILLER_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1924_ __dut__._2039_/B __dut__._2045_/B VGND VGND VPWR VPWR __dut__.__uuf__._1925_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1855_ __dut__.__uuf__._1877_/A __dut__.__uuf__._1855_/B __dut__.__uuf__._1855_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1856_/A sky130_fd_sc_hd__or3_4
XFILLER_138_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1786_ __dut__.__uuf__._1786_/A VGND VGND VPWR VPWR __dut__.__uuf__._1786_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_137_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1971_ __dut__._2213_/A __dut__._1971_/B VGND VGND VPWR VPWR __dut__._1971_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1336__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2407_ __dut__.__uuf__._2415_/CLK __dut__._2318_/X __dut__.__uuf__._1099_/X
+ VGND VGND VPWR VPWR __dut__._2319_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__212__A tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2338_ __dut__.__uuf__._2348_/CLK __dut__._2180_/X __dut__.__uuf__._1366_/X
+ VGND VGND VPWR VPWR __dut__._2181_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_121_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2523_ rst VGND VGND VPWR VPWR __dut__._2523_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2269_ __dut__.__uuf__._2270_/CLK __dut__._2042_/X __dut__.__uuf__._1608_/X
+ VGND VGND VPWR VPWR __dut__._2043_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_87_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2454_ rst VGND VGND VPWR VPWR __dut__._2454_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2385_ rst VGND VGND VPWR VPWR __dut__._2385_/Y sky130_fd_sc_hd__inv_2
X__dut__._1405_ __dut__._1433_/A __dut__._2656_/Q VGND VGND VPWR VPWR __dut__._1405_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_74_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1336_ __dut__._1282_/Y mc[21] __dut__._1335_/X VGND VGND VPWR VPWR __dut__._1336_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_215_ _292_/Q _290_/Q _231_/A VGND VGND VPWR VPWR _289_/D sky130_fd_sc_hd__o21a_4
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_146_ _308_/Q _237_/A VGND VGND VPWR VPWR _146_/X sky130_fd_sc_hd__and2_4
XFILLER_137_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_136_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2149__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_303_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1640_ __dut__.__uuf__._1642_/A VGND VGND VPWR VPWR __dut__.__uuf__._1640_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1571_ __dut__.__uuf__._1577_/A VGND VGND VPWR VPWR __dut__.__uuf__._1571_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1413__A __dut__.__uuf__._1711_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2612__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2123_ VGND VGND VPWR VPWR __dut__.__uuf__._2123_/HI tie[68] sky130_fd_sc_hd__conb_1
XFILLER_69_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2054_ __dut__.__uuf__._2054_/A VGND VGND VPWR VPWR __dut__.__uuf__._2054_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_84_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2308__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_72_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2170_ __dut__._2180_/A1 __dut__._2170_/A2 __dut__._2169_/X VGND VGND VPWR
+ VPWR __dut__._2170_/X sky130_fd_sc_hd__a21o_4
XFILLER_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2059__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1907_ __dut__.__uuf__._1907_/A VGND VGND VPWR VPWR __dut__.__uuf__._1909_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1838_ __dut__._1292_/X VGND VGND VPWR VPWR __dut__.__uuf__._1842_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_138_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1769_ __dut__.__uuf__._1769_/A VGND VGND VPWR VPWR __dut__._1980_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_119_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1954_ __dut__._2228_/A1 __dut__._1954_/A2 __dut__._1953_/X VGND VGND VPWR
+ VPWR __dut__._1954_/X sky130_fd_sc_hd__a21o_4
XFILLER_134_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2522__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1885_ __dut__._2313_/A __dut__._1885_/B VGND VGND VPWR VPWR __dut__._1885_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_153_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2506_ rst VGND VGND VPWR VPWR __dut__._2506_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_8_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2437_ rst VGND VGND VPWR VPWR __dut__._2437_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2368_ rst VGND VGND VPWR VPWR __dut__._2368_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__269__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1319_ _234_/Y __dut__._2636_/Q VGND VGND VPWR VPWR __dut__._1319_/X sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_3_4_0___dut__.__uuf__.__clk_source___A clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2299_ __dut__._2313_/A __dut__._2299_/B VGND VGND VPWR VPWR __dut__._2299_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_15_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2845__CLK __dut__._2845_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1601__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_129_ _129_/A VGND VGND VPWR VPWR _312_/D sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2432__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_253_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2607__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1511__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1623_ __dut__.__uuf__._1624_/A VGND VGND VPWR VPWR __dut__.__uuf__._1623_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1554_ __dut__.__uuf__._1543_/X __dut__.__uuf__._1538_/X __dut__._2101_/B
+ __dut__.__uuf__._1548_/X __dut__.__uuf__._1553_/X VGND VGND VPWR VPWR __dut__._2100_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1485_ __dut__.__uuf__._1507_/A VGND VGND VPWR VPWR __dut__.__uuf__._1485_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1670_ __dut__._1670_/A1 tie[62] __dut__._1669_/X VGND VGND VPWR VPWR __dut__._2754_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2106_ VGND VGND VPWR VPWR __dut__.__uuf__._2106_/HI tie[51] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2037_ __dut__.__uuf__._2037_/A __dut__.__uuf__._2037_/B __dut__.__uuf__._2037_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2038_/A sky130_fd_sc_hd__or3_4
XFILLER_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2222_ __dut__._2228_/A1 __dut__._2222_/A2 __dut__._2221_/X VGND VGND VPWR
+ VPWR __dut__._2222_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2280__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_72_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2153_ __dut__._2153_/A __dut__._2153_/B VGND VGND VPWR VPWR __dut__._2153_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2084_ __dut__._2084_/A1 __dut__._2084_/A2 __dut__._2083_/X VGND VGND VPWR
+ VPWR __dut__._2084_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2517__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_37_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1937_ __dut__._2327_/A __dut__._2887_/Q VGND VGND VPWR VPWR __dut__._1937_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1868_ __dut__._1868_/A1 tie[161] __dut__._1867_/X VGND VGND VPWR VPWR __dut__._2853_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1702__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1799_ __dut__._2213_/A __dut__._2818_/Q VGND VGND VPWR VPWR __dut__._1799_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1331__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2427__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1270_ __dut__.__uuf__._1429_/A VGND VGND VPWR VPWR __dut__.__uuf__._1270_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_7 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1766_/A1 sky130_fd_sc_hd__buf_2
X__dut__._2840_ clkbuf_opt_2_tck/A __dut__._2840_/D __dut__._2412_/Y VGND VGND VPWR
+ VPWR __dut__._2840_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1606_ __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR __dut__.__uuf__._1611_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_135_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2771_ __dut__._2865_/CLK __dut__._2771_/D __dut__._2481_/Y VGND VGND VPWR
+ VPWR __dut__._2771_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1537_ __dut__.__uuf__._1537_/A VGND VGND VPWR VPWR __dut__.__uuf__._1537_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1722_ __dut__._1722_/A1 tie[88] __dut__._1721_/X VGND VGND VPWR VPWR __dut__._2780_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1468_ __dut__.__uuf__._1455_/X __dut__.__uuf__._1450_/X __dut__._2141_/B
+ __dut__.__uuf__._1462_/X __dut__.__uuf__._1467_/X VGND VGND VPWR VPWR __dut__._2140_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_134_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1653_ __dut__._1661_/A __dut__._2745_/Q VGND VGND VPWR VPWR __dut__._1653_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1399_ __dut__.__uuf__._1398_/Y __dut__.__uuf__._1388_/X __dut__.__uuf__._1389_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1399_/X sky130_fd_sc_hd__o21a_4
XFILLER_134_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1584_ __dut__._1584_/A1 tie[19] __dut__._1583_/X VGND VGND VPWR VPWR __dut__._2711_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2690__CLK clkbuf_5_2_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2205_ __dut__._2213_/A __dut__._2205_/B VGND VGND VPWR VPWR __dut__._2205_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2136_ __dut__._2136_/A1 __dut__._2136_/A2 __dut__._2135_/X VGND VGND VPWR
+ VPWR __dut__._2136_/X sky130_fd_sc_hd__a21o_4
XFILLER_40_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2067_ __dut__._2213_/A __dut__._2067_/B VGND VGND VPWR VPWR __dut__._2067_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2176__A1 __dut__._2176_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_216_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_191 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2244_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_180 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2276_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_14 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1872_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_25 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1802_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_47 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1394_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_36 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2046_/A1 sky130_fd_sc_hd__buf_2
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2371_ __dut__.__uuf__._2372_/CLK __dut__._2246_/X __dut__.__uuf__._1206_/X
+ VGND VGND VPWR VPWR __dut__._2247_/B sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_69 psn_inst_psn_buff_73/A VGND VGND VPWR VPWR __dut__._2182_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_58 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1960_/A1 sky130_fd_sc_hd__buf_2
XFILLER_132_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1322_ __dut__.__uuf__._1315_/X __dut__.__uuf__._1321_/X __dut__._2199_/B
+ __dut__.__uuf__._1315_/X VGND VGND VPWR VPWR __dut__._2198_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1253_ __dut__.__uuf__._1355_/A VGND VGND VPWR VPWR __dut__.__uuf__._1269_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_113_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2620__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_opt_0_tck_A clkbuf_opt_1_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1184_ __dut__.__uuf__._1190_/A VGND VGND VPWR VPWR __dut__.__uuf__._1184_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_64_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2067__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2823_ clkbuf_5_1_0_tck/X __dut__._2823_/D __dut__._2429_/Y VGND VGND VPWR
+ VPWR __dut__._2823_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2754_ __dut__._2767_/CLK __dut__._2754_/D __dut__._2498_/Y VGND VGND VPWR
+ VPWR __dut__._2754_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1705_ __dut__._1705_/A __dut__._2771_/Q VGND VGND VPWR VPWR __dut__._1705_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_150_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2530__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2685_ __dut__._2744_/CLK __dut__._2685_/D __dut__._2567_/Y VGND VGND VPWR
+ VPWR __dut__._2685_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1636_ __dut__._1658_/A1 tie[45] __dut__._1635_/X VGND VGND VPWR VPWR __dut__._2737_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1567_ __dut__._1611_/A __dut__._2702_/Q VGND VGND VPWR VPWR __dut__._1567_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1498_ __dut__._1616_/A1 __dut__._1496_/X __dut__._1497_/X VGND VGND VPWR
+ VPWR __dut__._2680_/D sky130_fd_sc_hd__a21o_4
XFILLER_18_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2119_ __dut__._2149_/A __dut__._2119_/B VGND VGND VPWR VPWR __dut__._2119_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1372__A2 mc[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2440__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_166_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_333_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1940_ __dut__.__uuf__._1940_/A VGND VGND VPWR VPWR __dut__.__uuf__._1942_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1871_ __dut__.__uuf__._1871_/A VGND VGND VPWR VPWR __dut__.__uuf__._1871_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_51_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2615__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2423_ __dut__.__uuf__._2426_/CLK __dut__._2350_/X __dut__.__uuf__._1049_/X
+ VGND VGND VPWR VPWR __dut__._2351_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2354_ __dut__.__uuf__._2355_/CLK __dut__._2212_/X __dut__.__uuf__._1280_/X
+ VGND VGND VPWR VPWR __dut__._2213_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1305_ __dut__.__uuf__._1323_/A VGND VGND VPWR VPWR __dut__.__uuf__._1305_/X
+ sky130_fd_sc_hd__buf_2
Xclkbuf_3_3_0___dut__.__uuf__.__clk_source__ clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_7_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_132_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2285_ __dut__.__uuf__._2288_/CLK __dut__._2074_/X __dut__.__uuf__._1589_/X
+ VGND VGND VPWR VPWR __dut__._2075_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_87_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2470_ rst VGND VGND VPWR VPWR __dut__._2470_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1236_ __dut__.__uuf__._1236_/A VGND VGND VPWR VPWR __dut__.__uuf__._1260_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1421_ __dut__._1433_/A __dut__._2659_/Q VGND VGND VPWR VPWR __dut__._1421_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1167_ __dut__.__uuf__._1162_/X __dut__.__uuf__._1159_/X __dut__._2275_/B
+ __dut__._2277_/B __dut__.__uuf__._1156_/X VGND VGND VPWR VPWR __dut__._2274_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1352_ __dut__._1282_/Y mc[25] __dut__._1351_/X VGND VGND VPWR VPWR __dut__._1352_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1098_ __dut__.__uuf__._1087_/X __dut__.__uuf__._1084_/X __dut__._2321_/B
+ __dut__._2323_/B __dut__.__uuf__._1097_/X VGND VGND VPWR VPWR __dut__._2320_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1283_ __dut__._2627_/Q _234_/Y VGND VGND VPWR VPWR __dut__._1283_/X sky130_fd_sc_hd__and2_4
XFILLER_27_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_300_ _193_/A _300_/D trst VGND VGND VPWR VPWR _300_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1326__A __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_231_ _231_/A _231_/B VGND VGND VPWR VPWR _302_/D sky130_fd_sc_hd__and2_4
XFILLER_156_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_162_ _284_/Q _171_/B VGND VGND VPWR VPWR _283_/D sky130_fd_sc_hd__or2_4
XANTENNA___dut__._2525__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2806_ clkbuf_opt_1_tck/A __dut__._2806_/D __dut__._2446_/Y VGND VGND VPWR
+ VPWR __dut__._2806_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2737_ __dut__._2744_/CLK __dut__._2737_/D __dut__._2515_/Y VGND VGND VPWR
+ VPWR __dut__._2737_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2668_ __dut__._2680_/CLK __dut__._2668_/D __dut__._2584_/Y VGND VGND VPWR
+ VPWR __dut__._2668_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1619_ __dut__._1661_/A __dut__._2728_/Q VGND VGND VPWR VPWR __dut__._1619_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2364__CLK __dut__.__uuf__._2402_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2599_ rst VGND VGND VPWR VPWR __dut__._2599_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2435__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_283_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2070_ VGND VGND VPWR VPWR __dut__.__uuf__._2070_/HI tie[15] sky130_fd_sc_hd__conb_1
XFILLER_84_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1923_ __dut__._1324_/X VGND VGND VPWR VPWR __dut__.__uuf__._1927_/B
+ sky130_fd_sc_hd__inv_2
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1854_ __dut__.__uuf__._1821_/X __dut__.__uuf__._1852_/B __dut__.__uuf__._1852_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1855_/C sky130_fd_sc_hd__o21a_4
XFILLER_138_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1785_ __dut__._1987_/B __dut__._1993_/B VGND VGND VPWR VPWR __dut__.__uuf__._1786_/A
+ sky130_fd_sc_hd__and2_4
X__dut__._1970_ __dut__._2078_/A1 __dut__._1970_/A2 __dut__._1969_/X VGND VGND VPWR
+ VPWR __dut__._1970_/X sky130_fd_sc_hd__a21o_4
XFILLER_153_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2237__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1336__A2 mc[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2406_ __dut__.__uuf__._2412_/CLK __dut__._2316_/X __dut__.__uuf__._1102_/X
+ VGND VGND VPWR VPWR __dut__._2317_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2337_ __dut__.__uuf__._2348_/CLK __dut__._2178_/X __dut__.__uuf__._1371_/X
+ VGND VGND VPWR VPWR __dut__._2179_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_114_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2522_ rst VGND VGND VPWR VPWR __dut__._2522_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2268_ __dut__.__uuf__._2270_/CLK __dut__._2040_/X __dut__.__uuf__._1609_/X
+ VGND VGND VPWR VPWR __dut__._2041_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_59_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1219_ __dut__.__uuf__._1207_/X __dut__.__uuf__._1218_/X __dut__._2239_/B
+ __dut__._2241_/B __dut__.__uuf__._1215_/X VGND VGND VPWR VPWR __dut__._2238_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._2199_ VGND VGND VPWR VPWR __dut__.__uuf__._2199_/HI tie[144] sky130_fd_sc_hd__conb_1
XFILLER_142_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2453_ rst VGND VGND VPWR VPWR __dut__._2453_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1404_ __dut__._1282_/Y mp[5] __dut__._1403_/X VGND VGND VPWR VPWR __dut__._1404_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._2384_ rst VGND VGND VPWR VPWR __dut__._2384_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1335_ _234_/Y __dut__._2640_/Q VGND VGND VPWR VPWR __dut__._1335_/X sky130_fd_sc_hd__and2_4
XFILLER_43_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ _224_/B VGND VGND VPWR VPWR _231_/A sky130_fd_sc_hd__buf_2
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_145_ _237_/A VGND VGND VPWR VPWR _145_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_5_0_tck clkbuf_5_5_0_tck/A VGND VGND VPWR VPWR clkbuf_5_5_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_129_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1570_ __dut__.__uuf__._1564_/X __dut__.__uuf__._1559_/X __dut__._2093_/B
+ __dut__.__uuf__._1462_/A __dut__.__uuf__._1569_/X VGND VGND VPWR VPWR __dut__._2092_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_135_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2122_ VGND VGND VPWR VPWR __dut__.__uuf__._2122_/HI tie[67] sky130_fd_sc_hd__conb_1
XFILLER_130_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2053_ done __dut__.__uuf__._2052_/Y __dut__._1524_/X VGND VGND VPWR
+ VPWR __dut__._1956_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_69_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1906_ __dut__.__uuf__._1906_/A __dut__.__uuf__._1906_/B __dut__.__uuf__._1906_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1907_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1837_ __dut__.__uuf__._1829_/A __dut__.__uuf__._1834_/B __dut__.__uuf__._1836_/X
+ VGND VGND VPWR VPWR __dut__._2002_/A2 sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._2075__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1768_ __dut__.__uuf__._1768_/A __dut__.__uuf__._1768_/B __dut__.__uuf__._1768_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1769_/A sky130_fd_sc_hd__or3_4
X__dut__._1953_ __dut__._1953_/A __dut__._2688_/Q VGND VGND VPWR VPWR __dut__._1953_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1699_ __dut__._2339_/B __dut__.__uuf__._1695_/X __dut__._2275_/B
+ __dut__.__uuf__._1696_/X VGND VGND VPWR VPWR prod[22] sky130_fd_sc_hd__o22a_4
X__dut__._1884_ __dut__._1884_/A1 tie[169] __dut__._1883_/X VGND VGND VPWR VPWR __dut__._2861_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_106_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2797__CLK _270_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1419__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2505_ rst VGND VGND VPWR VPWR __dut__._2505_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2436_ rst VGND VGND VPWR VPWR __dut__._2436_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2367_ rst VGND VGND VPWR VPWR __dut__._2367_/Y sky130_fd_sc_hd__inv_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1318_ __dut__._1318_/A1 __dut__._1316_/X __dut__._1317_/X VGND VGND VPWR
+ VPWR __dut__._2635_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2402__CLK __dut__.__uuf__._2402_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2298_ __dut__._2356_/A1 __dut__._2298_/A2 __dut__._2297_/X VGND VGND VPWR
+ VPWR __dut__._2298_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_128_ _120_/Y _230_/A _124_/X _127_/X VGND VGND VPWR VPWR _129_/A sky130_fd_sc_hd__a211o_4
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1484__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1999__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1622_ __dut__.__uuf__._1624_/A VGND VGND VPWR VPWR __dut__.__uuf__._1622_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2623__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1553_ __dut__._1412_/X __dut__.__uuf__._1544_/X __dut__._2103_/B
+ __dut__.__uuf__._1549_/X VGND VGND VPWR VPWR __dut__.__uuf__._1553_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1484_ __dut__.__uuf__._1548_/A VGND VGND VPWR VPWR __dut__.__uuf__._1484_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2105_ VGND VGND VPWR VPWR __dut__.__uuf__._2105_/HI tie[50] sky130_fd_sc_hd__conb_1
XFILLER_96_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2036_ __dut__.__uuf__._1742_/A __dut__.__uuf__._2034_/B __dut__.__uuf__._2034_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2037_/C sky130_fd_sc_hd__o21a_4
X__dut__._2221_ __dut__._2221_/A __dut__._2221_/B VGND VGND VPWR VPWR __dut__._2221_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2152_ __dut__._2152_/A1 __dut__._2152_/A2 __dut__._2151_/X VGND VGND VPWR
+ VPWR __dut__._2152_/X sky130_fd_sc_hd__a21o_4
X__dut__._2083_ __dut__._2213_/A __dut__._2083_/B VGND VGND VPWR VPWR __dut__._2083_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2533__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1936_ __dut__._2328_/A1 prod[25] __dut__._1935_/X VGND VGND VPWR VPWR __dut__._2887_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1950__A2 done VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1867_ __dut__._2213_/A __dut__._2852_/Q VGND VGND VPWR VPWR __dut__._1867_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1798_ __dut__._1798_/A1 tie[126] __dut__._1797_/X VGND VGND VPWR VPWR __dut__._2818_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2419_ rst VGND VGND VPWR VPWR __dut__._2419_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1244__A __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2443__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_196_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2618__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_8 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1884_/A1 sky130_fd_sc_hd__buf_2
XFILLER_50_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1605_ __dut__.__uuf__._1605_/A VGND VGND VPWR VPWR __dut__.__uuf__._1605_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1536_ __dut__.__uuf__._1522_/X __dut__.__uuf__._1517_/X __dut__._2109_/B
+ __dut__.__uuf__._1527_/X __dut__.__uuf__._1535_/X VGND VGND VPWR VPWR __dut__._2108_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1932__A2 prod[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2770_ __dut__._2865_/CLK __dut__._2770_/D __dut__._2482_/Y VGND VGND VPWR
+ VPWR __dut__._2770_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1721_ __dut__._1729_/A __dut__._2779_/Q VGND VGND VPWR VPWR __dut__._1721_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1467_ __dut__._1500_/X __dut__.__uuf__._1457_/X __dut__._2143_/B
+ __dut__.__uuf__._1463_/X VGND VGND VPWR VPWR __dut__.__uuf__._1467_/X sky130_fd_sc_hd__o22a_4
XFILLER_150_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1652_ __dut__._1658_/A1 tie[53] __dut__._1651_/X VGND VGND VPWR VPWR __dut__._2745_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1696__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1398_ __dut__._2171_/B VGND VGND VPWR VPWR __dut__.__uuf__._1398_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2835__CLK __dut__._2845_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1583_ __dut__._1611_/A __dut__._2710_/Q VGND VGND VPWR VPWR __dut__._1583_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_85_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1448__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2019_ __dut__.__uuf__._2012_/A __dut__.__uuf__._2017_/B __dut__.__uuf__._1998_/X
+ VGND VGND VPWR VPWR __dut__._2070_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_150_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2204_ __dut__._2204_/A1 __dut__._2204_/A2 __dut__._2203_/X VGND VGND VPWR
+ VPWR __dut__._2204_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2528__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2135_ __dut__._2149_/A __dut__._2135_/B VGND VGND VPWR VPWR __dut__._2135_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2066_ __dut__._2066_/A1 __dut__._2066_/A2 __dut__._2065_/X VGND VGND VPWR
+ VPWR __dut__._2066_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1919_ __dut__._2327_/A __dut__._2878_/Q VGND VGND VPWR VPWR __dut__._1919_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1607__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2438__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_209_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_111_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_170 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1910_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_181 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2272_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_145_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_192 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1950_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_129_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_15 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1870_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_26 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1800_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_37 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2054_/A1 sky130_fd_sc_hd__buf_2
XFILLER_144_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2370_ __dut__.__uuf__._2372_/CLK __dut__._2244_/X __dut__.__uuf__._1210_/X
+ VGND VGND VPWR VPWR __dut__._2245_/B sky130_fd_sc_hd__dfrtp_4
Xpsn_inst_psn_buff_48 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1390_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_59 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2202_/A1 sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2858__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1321_ __dut__.__uuf__._1320_/Y __dut__.__uuf__._1309_/X __dut__.__uuf__._1311_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1321_/X sky130_fd_sc_hd__o21a_4
XFILLER_132_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1252_ __dut__.__uuf__._1655_/A VGND VGND VPWR VPWR __dut__.__uuf__._1355_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_113_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1678__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1183_ __dut__.__uuf__._1177_/X __dut__.__uuf__._1174_/X __dut__._2263_/B
+ __dut__._2265_/B __dut__.__uuf__._1171_/X VGND VGND VPWR VPWR __dut__._2262_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1850__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2083__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2822_ clkbuf_5_1_0_tck/X __dut__._2822_/D __dut__._2430_/Y VGND VGND VPWR
+ VPWR __dut__._2822_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_145_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2753_ __dut__._2865_/CLK __dut__._2753_/D __dut__._2499_/Y VGND VGND VPWR
+ VPWR __dut__._2753_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1519_ __dut__.__uuf__._1501_/X __dut__.__uuf__._1517_/X __dut__._2117_/B
+ __dut__.__uuf__._1506_/X __dut__.__uuf__._1518_/X VGND VGND VPWR VPWR __dut__._2116_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_151_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1704_ __dut__._1726_/A1 tie[79] __dut__._1703_/X VGND VGND VPWR VPWR __dut__._2771_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_77_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2684_ __dut__._2744_/CLK __dut__._2684_/D __dut__._2568_/Y VGND VGND VPWR
+ VPWR __dut__._2684_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1427__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1635_ __dut__._1661_/A __dut__._2736_/Q VGND VGND VPWR VPWR __dut__._1635_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_97_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1566_ __dut__._1566_/A1 tie[10] __dut__._1565_/X VGND VGND VPWR VPWR __dut__._2702_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_57_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1497_ __dut__._1617_/A __dut__._2679_/Q VGND VGND VPWR VPWR __dut__._1497_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2118_ __dut__._2118_/A1 __dut__._2118_/A2 __dut__._2117_/X VGND VGND VPWR
+ VPWR __dut__._2118_/X sky130_fd_sc_hd__a21o_4
XFILLER_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2049_ __dut__._2051_/A __dut__._2049_/B VGND VGND VPWR VPWR __dut__._2049_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1522__A __dut__.__uuf__._1564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2293__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_127_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_159_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1832__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_326_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1870_ __dut__._2019_/B __dut__._2025_/B VGND VGND VPWR VPWR __dut__.__uuf__._1871_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_149_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2422_ __dut__.__uuf__._2422_/CLK __dut__._2348_/X __dut__.__uuf__._1053_/X
+ VGND VGND VPWR VPWR __dut__._2349_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2353_ __dut__.__uuf__._2355_/CLK __dut__._2210_/X __dut__.__uuf__._1285_/X
+ VGND VGND VPWR VPWR __dut__._2211_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1304_ __dut__.__uuf__._1298_/X __dut__.__uuf__._1303_/X __dut__._2205_/B
+ __dut__.__uuf__._1298_/X VGND VGND VPWR VPWR __dut__._2204_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2284_ __dut__.__uuf__._2288_/CLK __dut__._2072_/X __dut__.__uuf__._1590_/X
+ VGND VGND VPWR VPWR __dut__._2073_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_115_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1235_ __dut__.__uuf__._1263_/A __dut__.__uuf__._1263_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1236_/A sky130_fd_sc_hd__or2_4
XFILLER_140_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1420_ __dut__._1282_/Y mp[8] __dut__._1419_/X VGND VGND VPWR VPWR __dut__._1420_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_28_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1166_ __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR __dut__.__uuf__._1166_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1351_ _234_/Y __dut__._2644_/Q VGND VGND VPWR VPWR __dut__._1351_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1097_ __dut__.__uuf__._1141_/A VGND VGND VPWR VPWR __dut__.__uuf__._1097_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1282_ _234_/Y VGND VGND VPWR VPWR __dut__._1282_/Y sky130_fd_sc_hd__inv_8
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_230_ _230_/A _296_/Q _303_/Q VGND VGND VPWR VPWR _231_/B sky130_fd_sc_hd__or3_4
XFILLER_23_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1999_ __dut__.__uuf__._1991_/A __dut__.__uuf__._1996_/B __dut__.__uuf__._1998_/X
+ VGND VGND VPWR VPWR __dut__._2062_/A2 sky130_fd_sc_hd__o21a_4
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_161_ _285_/Q _163_/B VGND VGND VPWR VPWR _284_/D sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_12_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._2805_ clkbuf_opt_1_tck/A __dut__._2805_/D __dut__._2447_/Y VGND VGND VPWR
+ VPWR __dut__._2805_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2541__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2736_ __dut__._2744_/CLK __dut__._2736_/D __dut__._2516_/Y VGND VGND VPWR
+ VPWR __dut__._2736_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2667_ __dut__._2726_/CLK __dut__._2667_/D __dut__._2585_/Y VGND VGND VPWR
+ VPWR __dut__._2667_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__302__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1618_ __dut__._1658_/A1 tie[36] __dut__._1617_/X VGND VGND VPWR VPWR __dut__._2728_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_65_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2598_ rst VGND VGND VPWR VPWR __dut__._2598_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1549_ __dut__._1549_/A __dut__._2693_/Q VGND VGND VPWR VPWR __dut__._1549_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1814__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1252__A __dut__.__uuf__._1655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2451__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_276_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1922_ __dut__.__uuf__._1915_/A __dut__.__uuf__._1920_/B __dut__.__uuf__._1890_/X
+ VGND VGND VPWR VPWR __dut__._2034_/A2 sky130_fd_sc_hd__o21a_4
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1853_ __dut__.__uuf__._1853_/A VGND VGND VPWR VPWR __dut__.__uuf__._1855_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2626__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2230__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1162__A __dut__.__uuf__._1177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1784_ __dut__._1532_/X VGND VGND VPWR VPWR __dut__.__uuf__._1788_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_138_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2405_ __dut__.__uuf__._2415_/CLK __dut__._2314_/X __dut__.__uuf__._1106_/X
+ VGND VGND VPWR VPWR __dut__._2315_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_145_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2361__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2336_ __dut__.__uuf__._2348_/CLK __dut__._2176_/X __dut__.__uuf__._1375_/X
+ VGND VGND VPWR VPWR __dut__._2177_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_126_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2521_ rst VGND VGND VPWR VPWR __dut__._2521_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2267_ __dut__.__uuf__._2270_/CLK __dut__._2038_/X __dut__.__uuf__._1610_/X
+ VGND VGND VPWR VPWR __dut__._2039_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2452_ rst VGND VGND VPWR VPWR __dut__._2452_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1218_ __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR __dut__.__uuf__._1218_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2198_ VGND VGND VPWR VPWR __dut__.__uuf__._2198_/HI tie[143] sky130_fd_sc_hd__conb_1
XFILLER_87_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1403_ _234_/Y __dut__._2657_/Q VGND VGND VPWR VPWR __dut__._1403_/X sky130_fd_sc_hd__and2_4
XFILLER_142_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2383_ rst VGND VGND VPWR VPWR __dut__._2383_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1149_ __dut__.__uuf__._1149_/A VGND VGND VPWR VPWR __dut__.__uuf__._1161_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1334_ __dut__._1346_/A1 __dut__._1332_/X __dut__._1333_/X VGND VGND VPWR
+ VPWR __dut__._2639_/D sky130_fd_sc_hd__a21o_4
XFILLER_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2536__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_213_ _229_/A _213_/B VGND VGND VPWR VPWR _224_/B sky130_fd_sc_hd__nor2_4
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_144_ _237_/A _141_/Y tdi _308_/Q _143_/Y VGND VGND VPWR VPWR _308_/D sky130_fd_sc_hd__a32o_4
XFILLER_143_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2719_ __dut__._2721_/CLK __dut__._2719_/D __dut__._2533_/Y VGND VGND VPWR
+ VPWR __dut__._2719_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2288__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_4_0_tck_A clkbuf_3_5_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2446__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__295__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2121_ VGND VGND VPWR VPWR __dut__.__uuf__._2121_/HI tie[66] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2052_ __dut__.__uuf__._2052_/A VGND VGND VPWR VPWR __dut__.__uuf__._2052_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_111_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1905_ __dut__._2031_/B __dut__._2037_/B __dut__.__uuf__._1904_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1906_/C sky130_fd_sc_hd__o21ai_4
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1836_ __dut__.__uuf__._1890_/A VGND VGND VPWR VPWR __dut__.__uuf__._1836_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1767_ __dut__.__uuf__._1766_/X __dut__.__uuf__._1763_/B __dut__.__uuf__._1763_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1768_/C sky130_fd_sc_hd__o21a_4
XANTENNA___dut__.__uuf__._2354__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_125_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1952_ __dut__._1952_/A1 tie[0] __dut__._1951_/X VGND VGND VPWR VPWR __dut__._2895_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1698_ __dut__._2337_/B __dut__.__uuf__._1695_/X __dut__._2273_/B
+ __dut__.__uuf__._1696_/X VGND VGND VPWR VPWR prod[21] sky130_fd_sc_hd__o22a_4
X__dut__._1883_ __dut__._2213_/A __dut__._2860_/Q VGND VGND VPWR VPWR __dut__._1883_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_119_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2319_ __dut__.__uuf__._2319_/CLK __dut__._2142_/X __dut__.__uuf__._1460_/X
+ VGND VGND VPWR VPWR __dut__._2143_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_75_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2504_ rst VGND VGND VPWR VPWR __dut__._2504_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1435__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2435_ rst VGND VGND VPWR VPWR __dut__._2435_/Y sky130_fd_sc_hd__inv_2
X__dut__._2366_ rst VGND VGND VPWR VPWR __dut__._2366_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1317_ __dut__._1325_/A __dut__._2634_/Q VGND VGND VPWR VPWR __dut__._1317_/X
+ sky130_fd_sc_hd__and2_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2297_ __dut__._2313_/A __dut__._2297_/B VGND VGND VPWR VPWR __dut__._2297_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_102_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_127_ _213_/B VGND VGND VPWR VPWR _127_/X sky130_fd_sc_hd__buf_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_141_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1484__A2 mp[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2227__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_81_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_239_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1621_ __dut__.__uuf__._1624_/A VGND VGND VPWR VPWR __dut__.__uuf__._1621_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_107_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1552_ __dut__.__uuf__._1558_/A VGND VGND VPWR VPWR __dut__.__uuf__._1552_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1483_ __dut__.__uuf__._1494_/A VGND VGND VPWR VPWR __dut__.__uuf__._1483_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2104_ VGND VGND VPWR VPWR __dut__.__uuf__._2104_/HI tie[49] sky130_fd_sc_hd__conb_1
XFILLER_57_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2035_ __dut__.__uuf__._2035_/A VGND VGND VPWR VPWR __dut__.__uuf__._2037_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._2220_ __dut__._2228_/A1 __dut__._2220_/A2 __dut__._2219_/X VGND VGND VPWR
+ VPWR __dut__._2220_/X sky130_fd_sc_hd__a21o_4
X__dut__._2151_ __dut__._2213_/A __dut__._2151_/B VGND VGND VPWR VPWR __dut__._2151_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2082_ __dut__._2082_/A1 __dut__._2082_/A2 __dut__._2081_/X VGND VGND VPWR
+ VPWR __dut__._2082_/X sky130_fd_sc_hd__a21o_4
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1819_ __dut__.__uuf__._1852_/A __dut__.__uuf__._1819_/B __dut__.__uuf__._1819_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1820_/A sky130_fd_sc_hd__or3_4
XANTENNA__234__A _304_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1935_ __dut__._2327_/A __dut__._2886_/Q VGND VGND VPWR VPWR __dut__._1935_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_153_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_4_0_tck clkbuf_5_5_0_tck/A VGND VGND VPWR VPWR clkbuf_5_4_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1866_ __dut__._1866_/A1 tie[160] __dut__._1865_/X VGND VGND VPWR VPWR __dut__._2852_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_79_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1797_ __dut__._2213_/A __dut__._2817_/Q VGND VGND VPWR VPWR __dut__._1797_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2418_ rst VGND VGND VPWR VPWR __dut__._2418_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2349_ __dut__._2349_/A __dut__._2349_/B VGND VGND VPWR VPWR __dut__._2349_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_16_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_330 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2147_/A
+ sky130_fd_sc_hd__buf_2
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_189_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1803__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1_0_tck_A clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_9 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1882_/A1 sky130_fd_sc_hd__buf_2
XFILLER_148_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1604_ __dut__.__uuf__._1605_/A VGND VGND VPWR VPWR __dut__.__uuf__._1604_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1535_ __dut__._1432_/X __dut__.__uuf__._1523_/X __dut__._2111_/B
+ __dut__.__uuf__._1528_/X VGND VGND VPWR VPWR __dut__.__uuf__._1535_/X sky130_fd_sc_hd__o22a_4
XFILLER_151_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1720_ __dut__._1722_/A1 tie[87] __dut__._1719_/X VGND VGND VPWR VPWR __dut__._2779_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_2_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1466_ __dut__.__uuf__._1472_/A VGND VGND VPWR VPWR __dut__.__uuf__._1466_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1651_ __dut__._1661_/A __dut__._2744_/Q VGND VGND VPWR VPWR __dut__._1651_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1397_ __dut__.__uuf__._1401_/A VGND VGND VPWR VPWR __dut__.__uuf__._1397_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_89_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1582_ __dut__._1584_/A1 tie[18] __dut__._1581_/X VGND VGND VPWR VPWR __dut__._2710_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1448__A2 mp[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2018_ __dut__.__uuf__._2018_/A VGND VGND VPWR VPWR __dut__._2072_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_85_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2203_ __dut__._2213_/A __dut__._2203_/B VGND VGND VPWR VPWR __dut__._2203_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_60_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2134_ __dut__._2136_/A1 __dut__._2134_/A2 __dut__._2133_/X VGND VGND VPWR
+ VPWR __dut__._2134_/X sky130_fd_sc_hd__a21o_4
XFILLER_26_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_42_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2065_ __dut__._2213_/A __dut__._2065_/B VGND VGND VPWR VPWR __dut__._2065_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2544__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1080__A __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1384__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1918_ __dut__._2328_/A1 prod[16] __dut__._1917_/X VGND VGND VPWR VPWR __dut__._2878_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1849_ __dut__._1853_/A __dut__._2843_/Q VGND VGND VPWR VPWR __dut__._1849_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2454__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpsn_inst_psn_buff_171 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2258_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_160 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1892_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA_psn_inst_psn_buff_104_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_182 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2274_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_193 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1658_/A1
+ sky130_fd_sc_hd__buf_4
XFILLER_145_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_16 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1868_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_38 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2056_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_27 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1798_/A1 sky130_fd_sc_hd__buf_2
XFILLER_133_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_49 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2094_/A1 sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1320_ __dut__._2201_/B VGND VGND VPWR VPWR __dut__.__uuf__._1320_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_144_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1251_ __dut__.__uuf__._1229_/A __dut__.__uuf__._1250_/X __dut__.__uuf__._1241_/B
+ __dut__._2227_/B __dut__.__uuf__._1247_/X VGND VGND VPWR VPWR __dut__._2226_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_140_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1182_ __dut__.__uuf__._1190_/A VGND VGND VPWR VPWR __dut__.__uuf__._1182_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_113_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1165__A __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2364__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2802__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2821_ clkbuf_5_1_0_tck/X __dut__._2821_/D __dut__._2431_/Y VGND VGND VPWR
+ VPWR __dut__._2821_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2752_ __dut__._2894_/CLK __dut__._2752_/D __dut__._2500_/Y VGND VGND VPWR
+ VPWR __dut__._2752_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1518_ __dut__._1448_/X __dut__.__uuf__._1502_/X __dut__._2119_/B
+ __dut__.__uuf__._1507_/X VGND VGND VPWR VPWR __dut__.__uuf__._1518_/X sky130_fd_sc_hd__o22a_4
XFILLER_145_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1703_ __dut__._1703_/A __dut__._2770_/Q VGND VGND VPWR VPWR __dut__._1703_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1449_ __dut__.__uuf__._1449_/A VGND VGND VPWR VPWR __dut__.__uuf__._1449_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2683_ __dut__._2744_/CLK __dut__._2683_/D __dut__._2569_/Y VGND VGND VPWR
+ VPWR __dut__._2683_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1634_ __dut__._1658_/A1 tie[44] __dut__._1633_/X VGND VGND VPWR VPWR __dut__._2736_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1565_ __dut__._1611_/A __dut__._2701_/Q VGND VGND VPWR VPWR __dut__._1565_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2539__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1496_ __dut__._1282_/Y mp[26] __dut__._1495_/X VGND VGND VPWR VPWR __dut__._1496_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1443__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2117_ __dut__._2149_/A __dut__._2117_/B VGND VGND VPWR VPWR __dut__._2117_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2048_ __dut__._2052_/A1 __dut__._2048_/A2 __dut__._2047_/X VGND VGND VPWR
+ VPWR __dut__._2048_/X sky130_fd_sc_hd__a21o_4
XFILLER_41_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2449__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_221_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_319_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2825__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1348__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2421_ __dut__.__uuf__._2422_/CLK __dut__._2346_/X __dut__.__uuf__._1057_/X
+ VGND VGND VPWR VPWR __dut__._2347_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_9_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2352_ __dut__.__uuf__._2355_/CLK __dut__._2208_/X __dut__.__uuf__._1291_/X
+ VGND VGND VPWR VPWR __dut__._2209_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1303_ __dut__.__uuf__._1302_/Y __dut__.__uuf__._2047_/A __dut__.__uuf__._1283_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1303_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._2283_ __dut__.__uuf__._2288_/CLK __dut__._2070_/X __dut__.__uuf__._1591_/X
+ VGND VGND VPWR VPWR __dut__._2071_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_99_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1234_ __dut__.__uuf__._1234_/A __dut__.__uuf__._1234_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1263_/B sky130_fd_sc_hd__or2_4
XFILLER_115_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1520__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1165_ __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR __dut__.__uuf__._1176_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1350_ __dut__._1354_/A1 __dut__._1348_/X __dut__._1349_/X VGND VGND VPWR
+ VPWR __dut__._2643_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1096_ __dut__.__uuf__._1102_/A VGND VGND VPWR VPWR __dut__.__uuf__._1096_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2359__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1281_ __dut__._2213_/A VGND VGND VPWR VPWR __dut__._1281_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1998_ __dut__.__uuf__._1998_/A VGND VGND VPWR VPWR __dut__.__uuf__._1998_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_156_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_160_ _286_/Q _171_/B VGND VGND VPWR VPWR _285_/D sky130_fd_sc_hd__or2_4
XFILLER_7_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2804_ clkbuf_5_5_0_tck/X __dut__._2804_/D __dut__._2448_/Y VGND VGND VPWR
+ VPWR __dut__._2804_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_156_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2735_ __dut__._2744_/CLK __dut__._2735_/D __dut__._2517_/Y VGND VGND VPWR
+ VPWR __dut__._2735_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2666_ __dut__._2726_/CLK __dut__._2666_/D __dut__._2586_/Y VGND VGND VPWR
+ VPWR __dut__._2666_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1617_ __dut__._1617_/A __dut__._2727_/Q VGND VGND VPWR VPWR __dut__._1617_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2597_ rst VGND VGND VPWR VPWR __dut__._2597_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1548_ __dut__._1548_/A1 tie[1] __dut__._1547_/X VGND VGND VPWR VPWR __dut__._2693_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_73_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1479_ _234_/Y __dut__._2676_/Q VGND VGND VPWR VPWR __dut__._1479_/X sky130_fd_sc_hd__and2_4
XFILLER_34_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2848__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_289_ _312_/CLK _289_/D trst VGND VGND VPWR VPWR _289_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_127_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0_tck_A clkbuf_3_1_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1750__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_171_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_269_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1921_ __dut__.__uuf__._1921_/A VGND VGND VPWR VPWR __dut__._2036_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1852_ __dut__.__uuf__._1852_/A __dut__.__uuf__._1852_/B __dut__.__uuf__._1852_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1853_/A sky130_fd_sc_hd__or3_4
XFILLER_60_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1783_ __dut__.__uuf__._1775_/A __dut__.__uuf__._1780_/B __dut__.__uuf__._1782_/X
+ VGND VGND VPWR VPWR __dut__._1982_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_20_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2404_ __dut__.__uuf__._2415_/CLK __dut__._2312_/X __dut__.__uuf__._1108_/X
+ VGND VGND VPWR VPWR __dut__._2313_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_126_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2335_ __dut__.__uuf__._2335_/CLK __dut__._2174_/X __dut__.__uuf__._1382_/X
+ VGND VGND VPWR VPWR __dut__._2175_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2520_ rst VGND VGND VPWR VPWR __dut__._2520_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2266_ __dut__.__uuf__._2270_/CLK __dut__._2036_/X __dut__.__uuf__._1611_/X
+ VGND VGND VPWR VPWR __dut__._2037_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2451_ rst VGND VGND VPWR VPWR __dut__._2451_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2197_ VGND VGND VPWR VPWR __dut__.__uuf__._2197_/HI tie[142] sky130_fd_sc_hd__conb_1
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1217_ __dut__.__uuf__._1220_/A VGND VGND VPWR VPWR __dut__.__uuf__._1217_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1402_ __dut__._1402_/A1 __dut__._1400_/X __dut__._1401_/X VGND VGND VPWR
+ VPWR __dut__._2656_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1148_ __dut__.__uuf__._1147_/X __dut__.__uuf__._1144_/X __dut__._2287_/B
+ __dut__._2289_/B __dut__.__uuf__._1141_/X VGND VGND VPWR VPWR __dut__._2286_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__.__uuf__._1618__A __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2283__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_142_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2382_ rst VGND VGND VPWR VPWR __dut__._2382_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1333_ __dut__._1341_/A __dut__._2637_/Q VGND VGND VPWR VPWR __dut__._1333_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1079_ __dut__.__uuf__._1086_/A VGND VGND VPWR VPWR __dut__.__uuf__._1079_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_70_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ tms VGND VGND VPWR VPWR _229_/A sky130_fd_sc_hd__inv_2
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_143_ _219_/A VGND VGND VPWR VPWR _143_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2552__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2718_ clkbuf_5_8_0_tck/X __dut__._2718_/D __dut__._2534_/Y VGND VGND VPWR
+ VPWR __dut__._2718_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2649_ clkbuf_5_3_0_tck/X __dut__._2649_/D __dut__._2603_/Y VGND VGND VPWR
+ VPWR __dut__._2649_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_38_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2462__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2120_ VGND VGND VPWR VPWR __dut__.__uuf__._2120_/HI tie[65] sky130_fd_sc_hd__conb_1
XFILLER_130_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2051_ __dut__.__uuf__._2051_/A __dut__._1957_/B __dut__.__uuf__._2051_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2052_/A sky130_fd_sc_hd__or3_4
XFILLER_96_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1904_ __dut__.__uuf__._1904_/A VGND VGND VPWR VPWR __dut__.__uuf__._1904_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1835_ __dut__.__uuf__._1835_/A VGND VGND VPWR VPWR __dut__._2004_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1766_ __dut__.__uuf__._2044_/A VGND VGND VPWR VPWR __dut__.__uuf__._1766_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_153_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2372__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1951_ __dut__._1951_/A __dut__._2894_/Q VGND VGND VPWR VPWR __dut__._1951_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1697_ __dut__._2335_/B __dut__.__uuf__._1695_/X __dut__._2271_/B
+ __dut__.__uuf__._1696_/X VGND VGND VPWR VPWR prod[20] sky130_fd_sc_hd__o22a_4
X__dut__._1882_ __dut__._1882_/A1 tie[168] __dut__._1881_/X VGND VGND VPWR VPWR __dut__._2860_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1714__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2318_ __dut__.__uuf__._2319_/CLK __dut__._2140_/X __dut__.__uuf__._1466_/X
+ VGND VGND VPWR VPWR __dut__._2141_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2503_ rst VGND VGND VPWR VPWR __dut__._2503_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2693__CLK clkbuf_5_2_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2249_ __dut__.__uuf__._2288_/CLK __dut__._2002_/X __dut__.__uuf__._1633_/X
+ VGND VGND VPWR VPWR __dut__._2003_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2434_ rst VGND VGND VPWR VPWR __dut__._2434_/Y sky130_fd_sc_hd__inv_2
X__dut__._2365_ rst VGND VGND VPWR VPWR __dut__._2365_/Y sky130_fd_sc_hd__inv_2
X__dut__._1316_ __dut__._1282_/Y mc[17] __dut__._1315_/X VGND VGND VPWR VPWR __dut__._1316_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2547__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1451__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2296_ __dut__._2356_/A1 __dut__._2296_/A2 __dut__._2295_/X VGND VGND VPWR
+ VPWR __dut__._2296_/X sky130_fd_sc_hd__a21o_4
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_126_ tms _255_/D _256_/Q _126_/D VGND VGND VPWR VPWR _213_/B sky130_fd_sc_hd__and4_4
XFILLER_98_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_134_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2457__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_301_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1620_ __dut__.__uuf__._1624_/A VGND VGND VPWR VPWR __dut__.__uuf__._1620_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1551_ __dut__.__uuf__._1543_/X __dut__.__uuf__._1538_/X __dut__._2103_/B
+ __dut__.__uuf__._1548_/X __dut__.__uuf__._1550_/X VGND VGND VPWR VPWR __dut__._2102_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1482_ __dut__.__uuf__._1478_/X __dut__.__uuf__._1473_/X __dut__._2135_/B
+ __dut__.__uuf__._1462_/X __dut__.__uuf__._1481_/X VGND VGND VPWR VPWR __dut__._2134_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2103_ VGND VGND VPWR VPWR __dut__.__uuf__._2103_/HI tie[48] sky130_fd_sc_hd__conb_1
XFILLER_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2034_ __dut__.__uuf__._2044_/A __dut__.__uuf__._2034_/B __dut__.__uuf__._2034_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2035_/A sky130_fd_sc_hd__or3_4
XFILLER_45_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2367__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2150_ __dut__._2150_/A1 __dut__._2150_/A2 __dut__._2149_/X VGND VGND VPWR
+ VPWR __dut__._2150_/X sky130_fd_sc_hd__a21o_4
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2321__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2081_ __dut__._2213_/A __dut__._2081_/B VGND VGND VPWR VPWR __dut__._2081_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_80_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1818_ __dut__._1999_/B __dut__._2005_/B __dut__.__uuf__._1817_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1819_/C sky130_fd_sc_hd__o21ai_4
XFILLER_40_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1749_ __dut__._1416_/X VGND VGND VPWR VPWR __dut__.__uuf__._1753_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_153_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1934_ __dut__._2328_/A1 prod[24] __dut__._1933_/X VGND VGND VPWR VPWR __dut__._2886_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1865_ __dut__._2213_/A __dut__._2851_/Q VGND VGND VPWR VPWR __dut__._1865_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1796_ __dut__._1796_/A1 tie[125] __dut__._1795_/X VGND VGND VPWR VPWR __dut__._2817_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_121_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_6_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2417_ rst VGND VGND VPWR VPWR __dut__._2417_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2348_ __dut__._2356_/A1 __dut__._2348_/A2 __dut__._2347_/X VGND VGND VPWR
+ VPWR __dut__._2348_/X sky130_fd_sc_hd__a21o_4
XFILLER_73_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2279_ __dut__._2279_/A __dut__._2279_/B VGND VGND VPWR VPWR __dut__._2279_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_320 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1341_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_331 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2215_/A
+ sky130_fd_sc_hd__buf_2
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_251_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1603_ __dut__.__uuf__._1605_/A VGND VGND VPWR VPWR __dut__.__uuf__._1603_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1534_ __dut__.__uuf__._1537_/A VGND VGND VPWR VPWR __dut__.__uuf__._1534_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1465_ __dut__.__uuf__._1455_/X __dut__.__uuf__._1450_/X __dut__._2143_/B
+ __dut__.__uuf__._1462_/X __dut__.__uuf__._1464_/X VGND VGND VPWR VPWR __dut__._2142_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1650_ __dut__._1658_/A1 tie[52] __dut__._1649_/X VGND VGND VPWR VPWR __dut__._2744_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1396_ __dut__.__uuf__._1393_/X __dut__.__uuf__._1395_/X __dut__._2171_/B
+ __dut__.__uuf__._1393_/X VGND VGND VPWR VPWR __dut__._2170_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1581_ __dut__._1611_/A __dut__._2709_/Q VGND VGND VPWR VPWR __dut__._1581_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2017_ __dut__.__uuf__._2037_/A __dut__.__uuf__._2017_/B __dut__.__uuf__._2017_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2018_/A sky130_fd_sc_hd__or3_4
XFILLER_85_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_6_0___dut__.__uuf__.__clk_source__ clkbuf_4_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2355_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_150_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2202_ __dut__._2202_/A1 __dut__._2202_/A2 __dut__._2201_/X VGND VGND VPWR
+ VPWR __dut__._2202_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._1268__B2 __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2133_ __dut__._2149_/A __dut__._2133_/B VGND VGND VPWR VPWR __dut__._2133_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_35_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2064_ __dut__._2064_/A1 __dut__._2064_/A2 __dut__._2063_/X VGND VGND VPWR
+ VPWR __dut__._2064_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1384__A2 mp[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1917_ __dut__._2327_/A __dut__._2877_/Q VGND VGND VPWR VPWR __dut__._1917_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2560__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1848_ __dut__._1854_/A1 tie[151] __dut__._1847_/X VGND VGND VPWR VPWR __dut__._2843_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1779_ __dut__._2213_/A __dut__._2808_/Q VGND VGND VPWR VPWR __dut__._1779_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_110_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_172 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2260_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_150 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1666_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_161 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1726_/A1
+ sky130_fd_sc_hd__buf_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_183 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2342_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_194 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2078_/A1 sky130_fd_sc_hd__buf_2
XFILLER_145_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_17 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1866_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_28 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1796_/A1 sky130_fd_sc_hd__buf_2
XANTENNA_psn_inst_psn_buff_299_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_39 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2060_/A1 sky130_fd_sc_hd__buf_2
XFILLER_144_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2470__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1250_ __dut__._2227_/B __dut__.__uuf__._1255_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1250_/X sky130_fd_sc_hd__or2_4
X__dut__.__uuf__._1181_ __dut__.__uuf__._1177_/X __dut__.__uuf__._1174_/X __dut__._2265_/B
+ __dut__._2267_/B __dut__.__uuf__._1171_/X VGND VGND VPWR VPWR __dut__._2264_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_140_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_3_0_tck clkbuf_5_3_0_tck/A VGND VGND VPWR VPWR clkbuf_5_3_0_tck/X sky130_fd_sc_hd__clkbuf_1
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._2820_ clkbuf_5_1_0_tck/X __dut__._2820_/D __dut__._2432_/Y VGND VGND VPWR
+ VPWR __dut__._2820_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2380__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2751_ __dut__._2894_/CLK __dut__._2751_/D __dut__._2501_/Y VGND VGND VPWR
+ VPWR __dut__._2751_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1517_ __dut__.__uuf__._1578_/A VGND VGND VPWR VPWR __dut__.__uuf__._1517_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_145_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1702_ __dut__._1726_/A1 tie[78] __dut__._1701_/X VGND VGND VPWR VPWR __dut__._2770_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2682_ clkbuf_5_3_0_tck/X __dut__._2682_/D __dut__._2570_/Y VGND VGND VPWR
+ VPWR __dut__._2682_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1448_ __dut__.__uuf__._1270_/X __dut__.__uuf__._1447_/X __dut__._2149_/B
+ __dut__.__uuf__._1270_/X VGND VGND VPWR VPWR __dut__._2148_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1633_ __dut__._1661_/A __dut__._2735_/Q VGND VGND VPWR VPWR __dut__._1633_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1379_ __dut__.__uuf__._1367_/X __dut__.__uuf__._1377_/X __dut__._2177_/B
+ __dut__.__uuf__._1378_/X VGND VGND VPWR VPWR __dut__._2176_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1564_ __dut__._1564_/A1 tie[9] __dut__._1563_/X VGND VGND VPWR VPWR __dut__._2701_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1495_ _234_/Y __dut__._2680_/Q VGND VGND VPWR VPWR __dut__._1495_/X sky130_fd_sc_hd__and2_4
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2555__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2116_ __dut__._2118_/A1 __dut__._2116_/A2 __dut__._2115_/X VGND VGND VPWR
+ VPWR __dut__._2116_/X sky130_fd_sc_hd__a21o_4
XFILLER_26_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2047_ __dut__._2051_/A __dut__._2047_/B VGND VGND VPWR VPWR __dut__._2047_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2627__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2306__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__289__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2465__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_214_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1348__A2 mc[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2420_ __dut__.__uuf__._2422_/CLK __dut__._2344_/X __dut__.__uuf__._1061_/X
+ VGND VGND VPWR VPWR __dut__._2345_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_117_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1809__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2351_ __dut__.__uuf__._2355_/CLK __dut__._2206_/X __dut__.__uuf__._1295_/X
+ VGND VGND VPWR VPWR __dut__._2207_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_126_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1302_ __dut__._2207_/B VGND VGND VPWR VPWR __dut__.__uuf__._1302_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2282_ __dut__.__uuf__._2282_/CLK __dut__._2068_/X __dut__.__uuf__._1592_/X
+ VGND VGND VPWR VPWR __dut__._2069_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_114_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1233_ __dut__._2217_/B VGND VGND VPWR VPWR __dut__.__uuf__._1234_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_115_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1520__A2 mp[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1164_ __dut__.__uuf__._1655_/A VGND VGND VPWR VPWR __dut__.__uuf__._1223_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_55_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1095_ __dut__.__uuf__._1087_/X __dut__.__uuf__._1084_/X __dut__._2323_/B
+ __dut__._2325_/B __dut__.__uuf__._1081_/X VGND VGND VPWR VPWR __dut__._2322_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1280_ rst VGND VGND VPWR VPWR __dut__._1280_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1284__A1 mc[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2375__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1997_ __dut__.__uuf__._1997_/A VGND VGND VPWR VPWR __dut__._2064_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2803_ clkbuf_5_5_0_tck/X __dut__._2803_/D __dut__._2449_/Y VGND VGND VPWR
+ VPWR __dut__._2803_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2734_ __dut__._2744_/CLK __dut__._2734_/D __dut__._2518_/Y VGND VGND VPWR
+ VPWR __dut__._2734_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2665_ __dut__._2726_/CLK __dut__._2665_/D __dut__._2587_/Y VGND VGND VPWR
+ VPWR __dut__._2665_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2596_ rst VGND VGND VPWR VPWR __dut__._2596_/Y sky130_fd_sc_hd__inv_2
X__dut__._1616_ __dut__._1616_/A1 tie[35] __dut__._1615_/X VGND VGND VPWR VPWR __dut__._2727_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_77_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1547_ __dut__._1951_/A __dut__._2895_/Q VGND VGND VPWR VPWR __dut__._1547_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1478_ __dut__._1616_/A1 __dut__._1476_/X __dut__._1477_/X VGND VGND VPWR
+ VPWR __dut__._2675_/D sky130_fd_sc_hd__a21o_4
XFILLER_61_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__311__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_288_ _288_/CLK _288_/D VGND VGND VPWR VPWR _288_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_164_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_331_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1920_ __dut__.__uuf__._1931_/A __dut__.__uuf__._1920_/B __dut__.__uuf__._1920_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1921_/A sky130_fd_sc_hd__or3_4
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2195__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1851_ __dut__._2011_/B __dut__._2017_/B __dut__.__uuf__._1850_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1852_/C sky130_fd_sc_hd__o21ai_4
XANTENNA___dut__._1811__B __dut__._2824_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1782_ __dut__.__uuf__._1890_/A VGND VGND VPWR VPWR __dut__.__uuf__._1782_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_118_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1539__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2403_ __dut__.__uuf__._2415_/CLK __dut__._2310_/X __dut__.__uuf__._1110_/X
+ VGND VGND VPWR VPWR __dut__._2311_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2334_ __dut__.__uuf__._2335_/CLK __dut__._2172_/X __dut__.__uuf__._1386_/X
+ VGND VGND VPWR VPWR __dut__._2173_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_126_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2265_ __dut__.__uuf__._2270_/CLK __dut__._2034_/X __dut__.__uuf__._1613_/X
+ VGND VGND VPWR VPWR __dut__._2035_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2450_ rst VGND VGND VPWR VPWR __dut__._2450_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2196_ VGND VGND VPWR VPWR __dut__.__uuf__._2196_/HI tie[141] sky130_fd_sc_hd__conb_1
XFILLER_120_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1216_ __dut__.__uuf__._1207_/X __dut__.__uuf__._1204_/X __dut__._2241_/B
+ __dut__._2243_/B __dut__.__uuf__._1215_/X VGND VGND VPWR VPWR __dut__._2240_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1401_ __dut__._1433_/A __dut__._2655_/Q VGND VGND VPWR VPWR __dut__._1401_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1147_ __dut__.__uuf__._1177_/A VGND VGND VPWR VPWR __dut__.__uuf__._1147_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2381_ rst VGND VGND VPWR VPWR __dut__._2381_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1332_ __dut__._1282_/Y mc[20] __dut__._1331_/X VGND VGND VPWR VPWR __dut__._1332_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1078_ __dut__.__uuf__._1072_/X __dut__.__uuf__._1069_/X __dut__._2333_/B
+ __dut__._2335_/B __dut__.__uuf__._1066_/X VGND VGND VPWR VPWR __dut__._2332_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_83_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ _203_/Y _207_/X _210_/X _252_/Q _244_/Q VGND VGND VPWR VPWR tdo sky130_fd_sc_hd__a32o_4
XFILLER_11_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_142_ _293_/Q _294_/Q VGND VGND VPWR VPWR _219_/A sky130_fd_sc_hd__or2_4
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2717_ clkbuf_5_9_0_tck/X __dut__._2717_/D __dut__._2535_/Y VGND VGND VPWR
+ VPWR __dut__._2717_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2648_ __dut__._2654_/CLK __dut__._2648_/D __dut__._2604_/Y VGND VGND VPWR
+ VPWR __dut__._2648_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1496__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2579_ rst VGND VGND VPWR VPWR __dut__._2579_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2815__CLK clkbuf_5_0_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1420__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1359__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_281_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2050_ __dut__._1524_/X __dut__.__uuf__._2050_/B VGND VGND VPWR VPWR
+ __dut__._1954_/A2 sky130_fd_sc_hd__and2_4
XFILLER_111_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1903_ __dut__._2031_/B __dut__._2037_/B VGND VGND VPWR VPWR __dut__.__uuf__._1904_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_80_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1834_ __dut__.__uuf__._1877_/A __dut__.__uuf__._1834_/B __dut__.__uuf__._1834_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1835_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1765_ __dut__.__uuf__._1765_/A VGND VGND VPWR VPWR __dut__.__uuf__._2044_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1950_ __dut__._1950_/A1 done __dut__._1949_/X VGND VGND VPWR VPWR __dut__._2894_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_153_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1696_ __dut__._1528_/X VGND VGND VPWR VPWR __dut__.__uuf__._1696_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1881_ __dut__._2213_/A __dut__._2859_/Q VGND VGND VPWR VPWR __dut__._1881_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_146_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2250__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2838__CLK clkbuf_opt_2_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2317_ __dut__.__uuf__._2319_/CLK __dut__._2138_/X __dut__.__uuf__._1469_/X
+ VGND VGND VPWR VPWR __dut__._2139_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2502_ rst VGND VGND VPWR VPWR __dut__._2502_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2248_ __dut__.__uuf__._2288_/CLK __dut__._2000_/X __dut__.__uuf__._1634_/X
+ VGND VGND VPWR VPWR __dut__._2001_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_153_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2433_ rst VGND VGND VPWR VPWR __dut__._2433_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2179_ VGND VGND VPWR VPWR __dut__.__uuf__._2179_/HI tie[124] sky130_fd_sc_hd__conb_1
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2364_ rst VGND VGND VPWR VPWR __dut__._2364_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1315_ _234_/Y __dut__._2635_/Q VGND VGND VPWR VPWR __dut__._1315_/X sky130_fd_sc_hd__and2_4
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_65_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2295_ __dut__._2313_/A __dut__._2295_/B VGND VGND VPWR VPWR __dut__._2295_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2563__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_125_ _254_/D _256_/D VGND VGND VPWR VPWR _126_/D sky130_fd_sc_hd__and2_4
XFILLER_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_127_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2473__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1550_ __dut__._1420_/X __dut__.__uuf__._1544_/X __dut__._2105_/B
+ __dut__.__uuf__._1549_/X VGND VGND VPWR VPWR __dut__.__uuf__._1550_/X sky130_fd_sc_hd__o22a_4
XFILLER_147_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1944__A2 prod[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1481_ __dut__._1488_/X __dut__.__uuf__._1480_/X __dut__._2137_/B
+ __dut__.__uuf__._1463_/X VGND VGND VPWR VPWR __dut__.__uuf__._1481_/X sky130_fd_sc_hd__o22a_4
XFILLER_128_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2102_ VGND VGND VPWR VPWR __dut__.__uuf__._2102_/HI tie[47] sky130_fd_sc_hd__conb_1
XFILLER_131_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2033_ __dut__._2079_/B __dut__._2085_/B __dut__.__uuf__._2032_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._2034_/C sky130_fd_sc_hd__o21ai_4
XFILLER_38_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2080_ __dut__._2080_/A1 __dut__._2080_/A2 __dut__._2079_/X VGND VGND VPWR
+ VPWR __dut__._2080_/X sky130_fd_sc_hd__a21o_4
XFILLER_52_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1817_ __dut__.__uuf__._1817_/A VGND VGND VPWR VPWR __dut__.__uuf__._1817_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_138_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2383__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1748_ __dut__.__uuf__._1983_/A VGND VGND VPWR VPWR __dut__.__uuf__._1798_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1933_ __dut__._2327_/A __dut__._2885_/Q VGND VGND VPWR VPWR __dut__._1933_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1679_ __dut__._2311_/B __dut__.__uuf__._1674_/X __dut__._2247_/B
+ __dut__.__uuf__._1675_/X VGND VGND VPWR VPWR prod[8] sky130_fd_sc_hd__o22a_4
XANTENNA___dut__._2660__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1864_ __dut__._1864_/A1 tie[159] __dut__._1863_/X VGND VGND VPWR VPWR __dut__._2851_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1795_ __dut__._2213_/A __dut__._2816_/Q VGND VGND VPWR VPWR __dut__._1795_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2416_ rst VGND VGND VPWR VPWR __dut__._2416_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2558__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2347_ __dut__._2349_/A __dut__._2347_/B VGND VGND VPWR VPWR __dut__._2347_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2278_ __dut__._2356_/A1 __dut__._2278_/A2 __dut__._2277_/X VGND VGND VPWR
+ VPWR __dut__._2278_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_310 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1289_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_321 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2051_/A
+ sky130_fd_sc_hd__buf_4
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._2296__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_332 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2153_/A
+ sky130_fd_sc_hd__buf_2
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2293__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._2468__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1602_ __dut__.__uuf__._1605_/A VGND VGND VPWR VPWR __dut__.__uuf__._1602_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_148_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1533_ __dut__.__uuf__._1522_/X __dut__.__uuf__._1517_/X __dut__._2111_/B
+ __dut__.__uuf__._1527_/X __dut__.__uuf__._1532_/X VGND VGND VPWR VPWR __dut__._2110_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1464_ __dut__._1508_/X __dut__.__uuf__._1457_/X __dut__._2145_/B
+ __dut__.__uuf__._1463_/X VGND VGND VPWR VPWR __dut__.__uuf__._1464_/X sky130_fd_sc_hd__o22a_4
XFILLER_104_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1395_ __dut__.__uuf__._1394_/Y __dut__.__uuf__._1388_/X __dut__.__uuf__._1389_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1395_/X sky130_fd_sc_hd__o21a_4
XANTENNA___dut__.__uuf__._1179__A __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1580_ __dut__._1580_/A1 tie[17] __dut__._1579_/X VGND VGND VPWR VPWR __dut__._2709_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_58_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2016_ __dut__.__uuf__._1983_/X __dut__.__uuf__._2014_/B __dut__.__uuf__._2014_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2017_/C sky130_fd_sc_hd__o21a_4
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2378__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1282__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2201_ __dut__._2213_/A __dut__._2201_/B VGND VGND VPWR VPWR __dut__._2201_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_150_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2132_ __dut__._2136_/A1 __dut__._2132_/A2 __dut__._2131_/X VGND VGND VPWR
+ VPWR __dut__._2132_/X sky130_fd_sc_hd__a21o_4
XFILLER_26_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2063_ __dut__._2213_/A __dut__._2063_/B VGND VGND VPWR VPWR __dut__._2063_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_28_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1916_ __dut__._2328_/A1 prod[15] __dut__._1915_/X VGND VGND VPWR VPWR __dut__._2877_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1457__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1847_ __dut__._1853_/A __dut__._2842_/Q VGND VGND VPWR VPWR __dut__._1847_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1778_ __dut__._1778_/A1 tie[116] __dut__._1777_/X VGND VGND VPWR VPWR __dut__._2808_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1844__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_140 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1616_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_173 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2262_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_151 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1668_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_162 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1894_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_195 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._2052_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_184 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2340_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_18 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1864_/A1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_29 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1794_/A1 sky130_fd_sc_hd__buf_2
XFILLER_145_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1367__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_194_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2311__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_152_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1180_ __dut__.__uuf__._1190_/A VGND VGND VPWR VPWR __dut__.__uuf__._1180_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_140_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1516_ __dut__.__uuf__._1516_/A VGND VGND VPWR VPWR __dut__.__uuf__._1516_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2750_ __dut__._2894_/CLK __dut__._2750_/D __dut__._2502_/Y VGND VGND VPWR
+ VPWR __dut__._2750_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2681_ __dut__._2744_/CLK __dut__._2681_/D __dut__._2571_/Y VGND VGND VPWR
+ VPWR __dut__._2681_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1701_ __dut__._1701_/A __dut__._2769_/Q VGND VGND VPWR VPWR __dut__._1701_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1447_ __dut__.__uuf__._1446_/Y __dut__.__uuf__._1438_/X __dut__.__uuf__._1337_/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._1447_/X sky130_fd_sc_hd__o21a_4
XFILLER_145_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1632_ __dut__._1658_/A1 tie[43] __dut__._1631_/X VGND VGND VPWR VPWR __dut__._2735_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1378_ __dut__.__uuf__._1393_/A VGND VGND VPWR VPWR __dut__.__uuf__._1378_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_77_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1563_ __dut__._1563_/A __dut__._2700_/Q VGND VGND VPWR VPWR __dut__._1563_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1826__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1494_ __dut__._1494_/A1 __dut__._1492_/X __dut__._1493_/X VGND VGND VPWR
+ VPWR __dut__._2679_/D sky130_fd_sc_hd__a21o_4
XFILLER_73_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2115_ __dut__._2149_/A __dut__._2115_/B VGND VGND VPWR VPWR __dut__._2115_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2046_ __dut__._2046_/A1 __dut__._2046_/A2 __dut__._2045_/X VGND VGND VPWR
+ VPWR __dut__._2046_/X sky130_fd_sc_hd__a21o_4
XFILLER_110_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2571__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2879_ __dut__._2892_/CLK __dut__._2879_/D __dut__._2373_/Y VGND VGND VPWR
+ VPWR __dut__._2879_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1915__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_19_0_tck clkbuf_4_9_0_tck/X VGND VGND VPWR VPWR __dut__._2865_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2481__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2350_ __dut__.__uuf__._2355_/CLK __dut__._2204_/X __dut__.__uuf__._1301_/X
+ VGND VGND VPWR VPWR __dut__._2205_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_132_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1301_ __dut__.__uuf__._1323_/A VGND VGND VPWR VPWR __dut__.__uuf__._1301_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2281_ __dut__.__uuf__._2288_/CLK __dut__._2066_/X __dut__.__uuf__._1593_/X
+ VGND VGND VPWR VPWR __dut__._2067_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_113_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1232_ __dut__._2221_/B VGND VGND VPWR VPWR __dut__.__uuf__._1263_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_141_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1825__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1163_ __dut__.__uuf__._1162_/X __dut__.__uuf__._1159_/X __dut__._2277_/B
+ __dut__._2279_/B __dut__.__uuf__._1156_/X VGND VGND VPWR VPWR __dut__._2276_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1094_ __dut__.__uuf__._1102_/A VGND VGND VPWR VPWR __dut__.__uuf__._1094_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1284__A2 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1192__A __dut__.__uuf__._1478_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1996_ __dut__.__uuf__._2037_/A __dut__.__uuf__._1996_/B __dut__.__uuf__._1996_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1997_/A sky130_fd_sc_hd__or3_4
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2391__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2802_ clkbuf_5_5_0_tck/X __dut__._2802_/D __dut__._2450_/Y VGND VGND VPWR
+ VPWR __dut__._2802_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2733_ __dut__._2744_/CLK __dut__._2733_/D __dut__._2519_/Y VGND VGND VPWR
+ VPWR __dut__._2733_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1735__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2664_ __dut__._2726_/CLK __dut__._2664_/D __dut__._2588_/Y VGND VGND VPWR
+ VPWR __dut__._2664_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2595_ rst VGND VGND VPWR VPWR __dut__._2595_/Y sky130_fd_sc_hd__inv_2
X__dut__._1615_ __dut__._1617_/A __dut__._2726_/Q VGND VGND VPWR VPWR __dut__._1615_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_95_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1546_ __dut__._1564_/A1 __dut__._1544_/X __dut__._1545_/X VGND VGND VPWR
+ VPWR __dut__._2692_/D sky130_fd_sc_hd__a21o_4
XFILLER_19_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1477_ __dut__._1477_/A __dut__._2674_/Q VGND VGND VPWR VPWR __dut__._1477_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2566__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2029_ __dut__._2029_/A __dut__._2029_/B VGND VGND VPWR VPWR __dut__._2029_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_155_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_287_ _288_/CLK _287_/D VGND VGND VPWR VPWR _287_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_2_0_tck clkbuf_5_3_0_tck/A VGND VGND VPWR VPWR clkbuf_5_2_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_157_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2476__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_324_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1850_ __dut__.__uuf__._1850_/A VGND VGND VPWR VPWR __dut__.__uuf__._1850_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1781_ __dut__.__uuf__._1781_/A VGND VGND VPWR VPWR __dut__._1984_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_137_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2402_ __dut__.__uuf__._2402_/CLK __dut__._2308_/X __dut__.__uuf__._1113_/X
+ VGND VGND VPWR VPWR __dut__._2309_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2333_ __dut__.__uuf__._2335_/CLK __dut__._2170_/X __dut__.__uuf__._1392_/X
+ VGND VGND VPWR VPWR __dut__._2171_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2264_ __dut__.__uuf__._2270_/CLK __dut__._2032_/X __dut__.__uuf__._1614_/X
+ VGND VGND VPWR VPWR __dut__._2033_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2195_ VGND VGND VPWR VPWR __dut__.__uuf__._2195_/HI tie[140] sky130_fd_sc_hd__conb_1
XFILLER_113_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._1215_ __dut__.__uuf__._1215_/A VGND VGND VPWR VPWR __dut__.__uuf__._1215_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2380_ rst VGND VGND VPWR VPWR __dut__._2380_/Y sky130_fd_sc_hd__inv_2
X__dut__._1400_ __dut__._1282_/Y mp[4] __dut__._1399_/X VGND VGND VPWR VPWR __dut__._1400_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1146_ __dut__.__uuf__._1146_/A VGND VGND VPWR VPWR __dut__.__uuf__._1146_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1331_ _234_/Y __dut__._2639_/Q VGND VGND VPWR VPWR __dut__._1331_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1077_ __dut__.__uuf__._1086_/A VGND VGND VPWR VPWR __dut__.__uuf__._1077_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2386__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_210_ _210_/A _210_/B VGND VGND VPWR VPWR _210_/X sky130_fd_sc_hd__or2_4
XFILLER_11_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1979_ __dut__.__uuf__._1979_/A VGND VGND VPWR VPWR __dut__.__uuf__._1979_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_141_ _294_/Q VGND VGND VPWR VPWR _141_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_psn_inst_psn_buff_10_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2716_ clkbuf_5_9_0_tck/X __dut__._2716_/D __dut__._2536_/Y VGND VGND VPWR
+ VPWR __dut__._2716_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2647_ __dut__._2654_/CLK __dut__._2647_/D __dut__._2605_/Y VGND VGND VPWR
+ VPWR __dut__._2647_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1496__A2 mp[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2578_ rst VGND VGND VPWR VPWR __dut__._2578_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1529_ __dut__._1529_/A __dut__._2687_/Q VGND VGND VPWR VPWR __dut__._1529_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_19_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1420__A2 mp[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_274_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1375__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1902_ __dut__._1316_/X VGND VGND VPWR VPWR __dut__.__uuf__._1906_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1833_ __dut__.__uuf__._1821_/X __dut__.__uuf__._1831_/B __dut__.__uuf__._1831_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1834_/C sky130_fd_sc_hd__o21a_4
XFILLER_40_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1764_ __dut__.__uuf__._1764_/A VGND VGND VPWR VPWR __dut__.__uuf__._1768_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_119_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1695_ __dut__.__uuf__._1702_/A VGND VGND VPWR VPWR __dut__.__uuf__._1695_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1880_ __dut__._1880_/A1 tie[167] __dut__._1879_/X VGND VGND VPWR VPWR __dut__._2859_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_118_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_9_0_tck clkbuf_4_9_0_tck/A VGND VGND VPWR VPWR clkbuf_4_9_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2316_ __dut__.__uuf__._2323_/CLK __dut__._2136_/X __dut__.__uuf__._1472_/X
+ VGND VGND VPWR VPWR __dut__._2137_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_121_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2501_ rst VGND VGND VPWR VPWR __dut__._2501_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1285__A tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2247_ __dut__.__uuf__._2288_/CLK __dut__._1998_/X __dut__.__uuf__._1635_/X
+ VGND VGND VPWR VPWR __dut__._1999_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2432_ rst VGND VGND VPWR VPWR __dut__._2432_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2178_ VGND VGND VPWR VPWR __dut__.__uuf__._2178_/HI tie[123] sky130_fd_sc_hd__conb_1
XFILLER_101_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2363_ rst VGND VGND VPWR VPWR __dut__._2363_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1129_ __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR __dut__.__uuf__._1188_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_90_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1314_ __dut__._1346_/A1 __dut__._1312_/X __dut__._1313_/X VGND VGND VPWR
+ VPWR __dut__._2634_/D sky130_fd_sc_hd__a21o_4
X__dut__._2294_ __dut__._2356_/A1 __dut__._2294_/A2 __dut__._2293_/X VGND VGND VPWR
+ VPWR __dut__._2294_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_58_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1380__A __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_124_ _235_/A _137_/B VGND VGND VPWR VPWR _124_/X sky130_fd_sc_hd__and2_4
XFILLER_152_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1923__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1480_ __dut__.__uuf__._1565_/A VGND VGND VPWR VPWR __dut__.__uuf__._1480_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2101_ VGND VGND VPWR VPWR __dut__.__uuf__._2101_/HI tie[46] sky130_fd_sc_hd__conb_1
XFILLER_69_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2032_ __dut__.__uuf__._2032_/A VGND VGND VPWR VPWR __dut__.__uuf__._2032_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_97_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1833__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1816_ __dut__._1999_/B __dut__._2005_/B VGND VGND VPWR VPWR __dut__.__uuf__._1817_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_148_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1396__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2805__CLK clkbuf_opt_1_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1747_ __dut__.__uuf__._1740_/A __dut__.__uuf__._1745_/B __dut__.__uuf__._1723_/X
+ VGND VGND VPWR VPWR __dut__._1970_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1932_ __dut__._2328_/A1 prod[23] __dut__._1931_/X VGND VGND VPWR VPWR __dut__._2885_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1678_ __dut__._2309_/B __dut__.__uuf__._1674_/X __dut__._2245_/B
+ __dut__.__uuf__._1675_/X VGND VGND VPWR VPWR prod[7] sky130_fd_sc_hd__o22a_4
XFILLER_134_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1863_ __dut__._2213_/A __dut__._2850_/Q VGND VGND VPWR VPWR __dut__._1863_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1794_ __dut__._1794_/A1 tie[124] __dut__._1793_/X VGND VGND VPWR VPWR __dut__._2816_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_121_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2415_ rst VGND VGND VPWR VPWR __dut__._2415_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1320__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2346_ __dut__._2356_/A1 __dut__._2346_/A2 __dut__._2345_/X VGND VGND VPWR
+ VPWR __dut__._2346_/X sky130_fd_sc_hd__a21o_4
X__dut__._2277_ __dut__._2277_/A __dut__._2277_/B VGND VGND VPWR VPWR __dut__._2277_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_311 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1545_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_300 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1505_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2574__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_322 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2095_/A
+ sky130_fd_sc_hd__buf_8
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_333 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2167_/A
+ sky130_fd_sc_hd__buf_2
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_237_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2240__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2484__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1601_ __dut__.__uuf__._1605_/A VGND VGND VPWR VPWR __dut__.__uuf__._1601_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_148_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1532_ __dut__._1436_/X __dut__.__uuf__._1523_/X __dut__._2113_/B
+ __dut__.__uuf__._1528_/X VGND VGND VPWR VPWR __dut__.__uuf__._1532_/X sky130_fd_sc_hd__o22a_4
XFILLER_116_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1463_ __dut__.__uuf__._1507_/A VGND VGND VPWR VPWR __dut__.__uuf__._1463_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_104_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1394_ __dut__._2173_/B VGND VGND VPWR VPWR __dut__.__uuf__._1394_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_103_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2015_ __dut__.__uuf__._2015_/A VGND VGND VPWR VPWR __dut__.__uuf__._2017_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2200_ __dut__._2200_/A1 __dut__._2200_/A2 __dut__._2199_/X VGND VGND VPWR
+ VPWR __dut__._2200_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2131_ __dut__._2149_/A __dut__._2131_/B VGND VGND VPWR VPWR __dut__._2131_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_26_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2394__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2062_ __dut__._2062_/A1 __dut__._2062_/A2 __dut__._2061_/X VGND VGND VPWR
+ VPWR __dut__._2062_/X sky130_fd_sc_hd__a21o_4
XFILLER_41_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1915_ __dut__._2327_/A __dut__._2876_/Q VGND VGND VPWR VPWR __dut__._1915_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_153_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2895_ clkbuf_5_0_0_tck/X __dut__._2895_/D __dut__._2626_/Y VGND VGND VPWR
+ VPWR __dut__._2895_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1846_ __dut__._1854_/A1 tie[150] __dut__._1845_/X VGND VGND VPWR VPWR __dut__._2842_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1777_ __dut__._2213_/A __dut__._2807_/Q VGND VGND VPWR VPWR __dut__._1777_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2569__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__305__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2329_ __dut__._2335_/A __dut__._2329_/B VGND VGND VPWR VPWR __dut__._2329_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_90_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_130 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1566_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_152 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1670_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_141 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1510_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_163 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1896_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_174 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2264_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_196 __dut__._1772_/A1 VGND VGND VPWR VPWR psn_inst_psn_buff_203/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_185 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2338_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_19 __dut__._1772_/A1 VGND VGND VPWR VPWR __dut__._1862_/A1 sky130_fd_sc_hd__buf_2
XFILLER_145_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_187_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1532__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2479__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1383__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1515_ __dut__.__uuf__._1501_/X __dut__.__uuf__._1495_/X __dut__._2119_/B
+ __dut__.__uuf__._1506_/X __dut__.__uuf__._1514_/X VGND VGND VPWR VPWR __dut__._2118_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_135_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2680_ __dut__._2680_/CLK __dut__._2680_/D __dut__._2572_/Y VGND VGND VPWR
+ VPWR __dut__._2680_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1700_ __dut__._1726_/A1 tie[77] __dut__._1699_/X VGND VGND VPWR VPWR __dut__._2769_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1446_ __dut__._2151_/B VGND VGND VPWR VPWR __dut__.__uuf__._1446_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_145_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1377_ __dut__.__uuf__._1376_/Y __dut__.__uuf__._1362_/X __dut__.__uuf__._1363_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1377_/X sky130_fd_sc_hd__o21a_4
X__dut__._1631_ __dut__._1661_/A __dut__._2734_/Q VGND VGND VPWR VPWR __dut__._1631_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2286__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1562_ __dut__._1564_/A1 tie[8] __dut__._1561_/X VGND VGND VPWR VPWR __dut__._2700_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2389__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1493_ __dut__._1493_/A __dut__._2678_/Q VGND VGND VPWR VPWR __dut__._1493_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2114_ __dut__._2118_/A1 __dut__._2114_/A2 __dut__._2113_/X VGND VGND VPWR
+ VPWR __dut__._2114_/X sky130_fd_sc_hd__a21o_4
XFILLER_26_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_40_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2045_ __dut__._2051_/A __dut__._2045_/B VGND VGND VPWR VPWR __dut__._2045_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1762__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2878_ __dut__._2892_/CLK __dut__._2878_/D __dut__._2374_/Y VGND VGND VPWR
+ VPWR __dut__._2878_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1829_ __dut__._1853_/A __dut__._2833_/Q VGND VGND VPWR VPWR __dut__._1829_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_79_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._2299__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1931__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_102_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__298__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2280_ __dut__.__uuf__._2288_/CLK __dut__._2064_/X __dut__.__uuf__._1595_/X
+ VGND VGND VPWR VPWR __dut__._2065_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1300_ __dut__.__uuf__._1355_/A VGND VGND VPWR VPWR __dut__.__uuf__._1323_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1231_ __dut__.__uuf__._1249_/A VGND VGND VPWR VPWR __dut__.__uuf__._1231_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_141_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1162_ __dut__.__uuf__._1177_/A VGND VGND VPWR VPWR __dut__.__uuf__._1162_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1093_ __dut__.__uuf__._1087_/X __dut__.__uuf__._1084_/X __dut__._2325_/B
+ __dut__._2327_/B __dut__.__uuf__._1081_/X VGND VGND VPWR VPWR __dut__._2324_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_28_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1841__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1473__A __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1995_ __dut__.__uuf__._1983_/X __dut__.__uuf__._1993_/B __dut__.__uuf__._1993_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1996_/C sky130_fd_sc_hd__o21a_4
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2801_ clkbuf_opt_2_tck/A __dut__._2801_/D __dut__._2451_/Y VGND VGND VPWR
+ VPWR __dut__._2801_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1744__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2732_ __dut__._2744_/CLK __dut__._2732_/D __dut__._2520_/Y VGND VGND VPWR
+ VPWR __dut__._2732_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2696__CLK clkbuf_5_2_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1429_ __dut__.__uuf__._1429_/A VGND VGND VPWR VPWR __dut__.__uuf__._1429_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_78_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2663_ __dut__._2726_/CLK __dut__._2663_/D __dut__._2589_/Y VGND VGND VPWR
+ VPWR __dut__._2663_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1614_ __dut__._1616_/A1 tie[34] __dut__._1613_/X VGND VGND VPWR VPWR __dut__._2726_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2594_ rst VGND VGND VPWR VPWR __dut__._2594_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1545_ __dut__._1545_/A __dut__._2691_/Q VGND VGND VPWR VPWR __dut__._1545_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_88_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1751__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1476_ __dut__._1282_/Y mp[21] __dut__._1475_/X VGND VGND VPWR VPWR __dut__._1476_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_73_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2301__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2028_ __dut__._2030_/A1 __dut__._2028_/A2 __dut__._2027_/X VGND VGND VPWR
+ VPWR __dut__._2028_/X sky130_fd_sc_hd__a21o_4
X_286_ _288_/CLK _286_/D VGND VGND VPWR VPWR _286_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._2582__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_317_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1780_ __dut__.__uuf__._1823_/A __dut__.__uuf__._1780_/B __dut__.__uuf__._1780_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1781_/A sky130_fd_sc_hd__or3_4
XANTENNA___dut__._2492__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1726__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2401_ __dut__.__uuf__._2402_/CLK __dut__._2306_/X __dut__.__uuf__._1116_/X
+ VGND VGND VPWR VPWR __dut__._2307_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2332_ __dut__.__uuf__._2335_/CLK __dut__._2168_/X __dut__.__uuf__._1397_/X
+ VGND VGND VPWR VPWR __dut__._2169_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2263_ __dut__.__uuf__._2270_/CLK __dut__._2030_/X __dut__.__uuf__._1615_/X
+ VGND VGND VPWR VPWR __dut__._2031_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2194_ VGND VGND VPWR VPWR __dut__.__uuf__._2194_/HI tie[139] sky130_fd_sc_hd__conb_1
XFILLER_87_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1214_ __dut__.__uuf__._1220_/A VGND VGND VPWR VPWR __dut__.__uuf__._1214_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_75_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1145_ __dut__.__uuf__._1133_/X __dut__.__uuf__._1144_/X __dut__._2289_/B
+ __dut__._2291_/B __dut__.__uuf__._1141_/X VGND VGND VPWR VPWR __dut__._2288_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1076_ __dut__.__uuf__._1072_/X __dut__.__uuf__._1069_/X __dut__._2335_/B
+ __dut__._2337_/B __dut__.__uuf__._1066_/X VGND VGND VPWR VPWR __dut__._2334_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1330_ __dut__._1330_/A1 __dut__._1328_/X __dut__._1329_/X VGND VGND VPWR
+ VPWR __dut__._2638_/D sky130_fd_sc_hd__a21o_4
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1571__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2324__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1978_ __dut__._2059_/B __dut__._2065_/B VGND VGND VPWR VPWR __dut__.__uuf__._1979_/A
+ sky130_fd_sc_hd__and2_4
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_140_ _293_/Q VGND VGND VPWR VPWR _237_/A sky130_fd_sc_hd__buf_2
XFILLER_51_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_18_0_tck clkbuf_4_9_0_tck/X VGND VGND VPWR VPWR __dut__._2767_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2715_ clkbuf_5_9_0_tck/X __dut__._2715_/D __dut__._2537_/Y VGND VGND VPWR
+ VPWR __dut__._2715_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2646_ __dut__._2654_/CLK __dut__._2646_/D __dut__._2606_/Y VGND VGND VPWR
+ VPWR __dut__._2646_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2577_ rst VGND VGND VPWR VPWR __dut__._2577_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2577__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1528_ __dut__._1282_/Y prod_sel __dut__._1527_/X VGND VGND VPWR VPWR __dut__._1528_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1459_ _234_/Y __dut__._2671_/Q VGND VGND VPWR VPWR __dut__._1459_/X sky130_fd_sc_hd__and2_4
XFILLER_34_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_269_ _271_/CLK _269_/D VGND VGND VPWR VPWR _269_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1708__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_267_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2487__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1391__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1901_ __dut__.__uuf__._1894_/A __dut__.__uuf__._1899_/B __dut__.__uuf__._1890_/X
+ VGND VGND VPWR VPWR __dut__._2026_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_52_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1832_ __dut__.__uuf__._1832_/A VGND VGND VPWR VPWR __dut__.__uuf__._1834_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_80_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1763_ __dut__.__uuf__._1798_/A __dut__.__uuf__._1763_/B __dut__.__uuf__._1763_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1764_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1694_ __dut__._2333_/B __dut__.__uuf__._1688_/X __dut__._2269_/B
+ __dut__.__uuf__._1689_/X VGND VGND VPWR VPWR prod[19] sky130_fd_sc_hd__o22a_4
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2315_ __dut__.__uuf__._2323_/CLK __dut__._2134_/X __dut__.__uuf__._1477_/X
+ VGND VGND VPWR VPWR __dut__._2135_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2500_ rst VGND VGND VPWR VPWR __dut__._2500_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1285__B __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2246_ __dut__.__uuf__._2288_/CLK __dut__._1996_/X __dut__.__uuf__._1636_/X
+ VGND VGND VPWR VPWR __dut__._1997_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2431_ rst VGND VGND VPWR VPWR __dut__._2431_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2177_ VGND VGND VPWR VPWR __dut__.__uuf__._2177_/HI tie[122] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2397__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2362_ rst VGND VGND VPWR VPWR __dut__._2362_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1128_ __dut__.__uuf__._1132_/A VGND VGND VPWR VPWR __dut__.__uuf__._1128_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1313_ __dut__._1313_/A __dut__._2633_/Q VGND VGND VPWR VPWR __dut__._1313_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2293_ __dut__._2313_/A __dut__._2293_/B VGND VGND VPWR VPWR __dut__._2293_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1059_ __dut__.__uuf__._1058_/X __dut__.__uuf__._1055_/X __dut__._2347_/B
+ __dut__._2349_/B __dut__.__uuf__._1051_/X VGND VGND VPWR VPWR __dut__._2346_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_71_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_1_0_tck clkbuf_5_1_0_tck/A VGND VGND VPWR VPWR clkbuf_5_1_0_tck/X sky130_fd_sc_hd__clkbuf_1
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1661__A __dut__.__uuf__._2054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_123_ _289_/Q VGND VGND VPWR VPWR _137_/B sky130_fd_sc_hd__inv_2
XFILLER_137_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2629_ __dut__._2357_/B __dut__._2629_/D __dut__._2623_/Y VGND VGND VPWR
+ VPWR __dut__._2629_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1836__A __dut__.__uuf__._1890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0___dut__.__uuf__.__clk_source__ clkbuf_2_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2354__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2100_ VGND VGND VPWR VPWR __dut__.__uuf__._2100_/HI tie[45] sky130_fd_sc_hd__conb_1
XFILLER_111_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2031_ __dut__._2079_/B __dut__._2085_/B VGND VGND VPWR VPWR __dut__.__uuf__._2032_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_97_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1815_ __dut__._1544_/X VGND VGND VPWR VPWR __dut__.__uuf__._1819_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1396__A2 mp[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1746_ __dut__.__uuf__._1746_/A VGND VGND VPWR VPWR __dut__._1972_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1931_ __dut__._2327_/A __dut__._2884_/Q VGND VGND VPWR VPWR __dut__._1931_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_5_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1677_ __dut__._2307_/B __dut__.__uuf__._1674_/X __dut__._2243_/B
+ __dut__.__uuf__._1675_/X VGND VGND VPWR VPWR prod[6] sky130_fd_sc_hd__o22a_4
XFILLER_134_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1862_ __dut__._1862_/A1 tie[158] __dut__._1861_/X VGND VGND VPWR VPWR __dut__._2850_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1793_ __dut__._1793_/A __dut__._2815_/Q VGND VGND VPWR VPWR __dut__._1793_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1856__B1 __dut__._1855_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._2229_ __dut__.__uuf__._2355_/CLK __dut__._1962_/X __dut__.__uuf__._1657_/X
+ VGND VGND VPWR VPWR __dut__._1963_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2414_ rst VGND VGND VPWR VPWR __dut__._2414_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1320__A2 mc[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2345_ __dut__._2349_/A __dut__._2345_/B VGND VGND VPWR VPWR __dut__._2345_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_56_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2276_ __dut__._2276_/A1 __dut__._2276_/A2 __dut__._2275_/X VGND VGND VPWR
+ VPWR __dut__._2276_/X sky130_fd_sc_hd__a21o_4
XFILLER_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_312 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2031_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_301 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1533_/A
+ sky130_fd_sc_hd__buf_2
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_323 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1433_/A
+ sky130_fd_sc_hd__buf_4
Xpsn_inst_psn_buff_334 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2213_/A
+ sky130_fd_sc_hd__buf_8
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2590__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0_tck clkbuf_4_9_0_tck/A VGND VGND VPWR VPWR clkbuf_4_8_0_tck/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_psn_inst_psn_buff_132_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1600_ __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR __dut__.__uuf__._1605_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_147_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1531_ __dut__.__uuf__._1537_/A VGND VGND VPWR VPWR __dut__.__uuf__._1531_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_144_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1462_ __dut__.__uuf__._1462_/A VGND VGND VPWR VPWR __dut__.__uuf__._1462_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2005__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1393_ __dut__.__uuf__._1393_/A VGND VGND VPWR VPWR __dut__.__uuf__._1393_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1838__B1 __dut__._1837_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1302__A2 __dut__._1300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2014_ __dut__.__uuf__._2014_/A __dut__.__uuf__._2014_/B __dut__.__uuf__._2014_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2015_/A sky130_fd_sc_hd__or3_4
XFILLER_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2130_ __dut__._2136_/A1 __dut__._2130_/A2 __dut__._2129_/X VGND VGND VPWR
+ VPWR __dut__._2130_/X sky130_fd_sc_hd__a21o_4
XFILLER_38_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2061_ __dut__._2213_/A __dut__._2061_/B VGND VGND VPWR VPWR __dut__._2061_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1729_ __dut__._1967_/B __dut__._1973_/B VGND VGND VPWR VPWR __dut__.__uuf__._1730_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_138_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1914_ __dut__._2328_/A1 prod[14] __dut__._1913_/X VGND VGND VPWR VPWR __dut__._2876_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_153_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2894_ __dut__._2894_/CLK __dut__._2894_/D __dut__._1280_/Y VGND VGND VPWR
+ VPWR __dut__._2894_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1845_ __dut__._1853_/A __dut__._2841_/Q VGND VGND VPWR VPWR __dut__._1845_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1776_ __dut__._1776_/A1 tie[115] __dut__._1775_/X VGND VGND VPWR VPWR __dut__._2807_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_4_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2585__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2328_ __dut__._2328_/A1 __dut__._2328_/A2 __dut__._2327_/X VGND VGND VPWR
+ VPWR __dut__._2328_/X sky130_fd_sc_hd__a21o_4
X__dut__._2259_ __dut__._2259_/A __dut__._2259_/B VGND VGND VPWR VPWR __dut__._2259_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_120 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2032_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_153 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1672_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_131 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1604_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_142 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1530_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_164 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1898_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_175 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2324_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_186 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1854_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_197 psn_inst_psn_buff_203/A VGND VGND VPWR VPWR __dut__._2062_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1929__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1532__A2 mc[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1296__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2495__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1839__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._1514_ __dut__._1452_/X __dut__.__uuf__._1502_/X __dut__._2121_/B
+ __dut__.__uuf__._1507_/X VGND VGND VPWR VPWR __dut__.__uuf__._1514_/X sky130_fd_sc_hd__o22a_4
XFILLER_135_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1445_ __dut__.__uuf__._1449_/A VGND VGND VPWR VPWR __dut__.__uuf__._1445_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1376_ __dut__._2179_/B VGND VGND VPWR VPWR __dut__.__uuf__._1376_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1630_ __dut__._1658_/A1 tie[42] __dut__._1629_/X VGND VGND VPWR VPWR __dut__._2734_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_131_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1561_ __dut__._1563_/A __dut__._2699_/Q VGND VGND VPWR VPWR __dut__._1561_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1492_ __dut__._1282_/Y mp[25] __dut__._1491_/X VGND VGND VPWR VPWR __dut__._1492_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2113_ __dut__._2149_/A __dut__._2113_/B VGND VGND VPWR VPWR __dut__._2113_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_26_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2044_ __dut__._2044_/A1 __dut__._2044_/A2 __dut__._2043_/X VGND VGND VPWR
+ VPWR __dut__._2044_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_33_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1749__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2877_ __dut__._2892_/CLK __dut__._2877_/D __dut__._2375_/Y VGND VGND VPWR
+ VPWR __dut__._2877_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1828_ __dut__._1854_/A1 tie[141] __dut__._1827_/X VGND VGND VPWR VPWR __dut__._2833_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2230__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2818__CLK clkbuf_5_0_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1759_ __dut__._1853_/A __dut__._2798_/Q VGND VGND VPWR VPWR __dut__._1759_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_96_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_297_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1230_ __dut__.__uuf__._1221_/X __dut__.__uuf__._1218_/X __dut__._2231_/B
+ __dut__._2233_/B __dut__.__uuf__._1229_/X VGND VGND VPWR VPWR __dut__._2230_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_113_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1161_ __dut__.__uuf__._1161_/A VGND VGND VPWR VPWR __dut__.__uuf__._1161_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_141_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1092_ __dut__.__uuf__._1102_/A VGND VGND VPWR VPWR __dut__.__uuf__._1092_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1994_ __dut__.__uuf__._1994_/A VGND VGND VPWR VPWR __dut__.__uuf__._1996_/B
+ sky130_fd_sc_hd__inv_2
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2053__A1 done VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2800_ clkbuf_opt_2_tck/A __dut__._2800_/D __dut__._2452_/Y VGND VGND VPWR
+ VPWR __dut__._2800_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._2731_ __dut__._2744_/CLK __dut__._2731_/D __dut__._2521_/Y VGND VGND VPWR
+ VPWR __dut__._2731_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2662_ __dut__._2726_/CLK __dut__._2662_/D __dut__._2590_/Y VGND VGND VPWR
+ VPWR __dut__._2662_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1428_ __dut__.__uuf__._1427_/Y __dut__.__uuf__._1413_/X __dut__.__uuf__._1414_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1428_/X sky130_fd_sc_hd__o21a_4
XFILLER_49_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1613_ __dut__._1617_/A __dut__._2725_/Q VGND VGND VPWR VPWR __dut__._1613_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2593_ rst VGND VGND VPWR VPWR __dut__._2593_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1359_ __dut__.__uuf__._1353_/X __dut__.__uuf__._1358_/X __dut__._2185_/B
+ __dut__.__uuf__._1353_/X VGND VGND VPWR VPWR __dut__._2184_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1544_ __dut__._1282_/Y mc[9] __dut__._1543_/X VGND VGND VPWR VPWR __dut__._1544_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1475_ _234_/Y __dut__._2675_/Q VGND VGND VPWR VPWR __dut__._1475_/X sky130_fd_sc_hd__and2_4
XFILLER_100_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_2_0___dut__.__uuf__.__clk_source__ clkbuf_4_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2319_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__.__uuf__._1664__A __dut__._1528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1680__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1432__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2027_ __dut__._2029_/A __dut__._2027_/B VGND VGND VPWR VPWR __dut__._2027_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_285_ _288_/CLK _285_/D VGND VGND VPWR VPWR _285_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1479__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_7_0___dut__.__uuf__.__clk_source___A clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_212_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2400_ __dut__.__uuf__._2402_/CLK __dut__._2304_/X __dut__.__uuf__._1121_/X
+ VGND VGND VPWR VPWR __dut__._2305_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_145_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2331_ __dut__.__uuf__._2335_/CLK __dut__._2166_/X __dut__.__uuf__._1401_/X
+ VGND VGND VPWR VPWR __dut__._2167_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2262_ __dut__.__uuf__._2270_/CLK __dut__._2028_/X __dut__.__uuf__._1616_/X
+ VGND VGND VPWR VPWR __dut__._2029_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1213_ __dut__.__uuf__._1207_/X __dut__.__uuf__._1204_/X __dut__._2243_/B
+ __dut__._2245_/B __dut__.__uuf__._1200_/X VGND VGND VPWR VPWR __dut__._2242_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._2193_ VGND VGND VPWR VPWR __dut__.__uuf__._2193_/HI tie[138] sky130_fd_sc_hd__conb_1
XFILLER_102_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2013__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1144_ __dut__.__uuf__._1188_/A VGND VGND VPWR VPWR __dut__.__uuf__._1144_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1075_ __dut__.__uuf__._1086_/A VGND VGND VPWR VPWR __dut__.__uuf__._1075_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_28_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1977_ __dut__._1348_/X VGND VGND VPWR VPWR __dut__.__uuf__._1981_/B
+ sky130_fd_sc_hd__inv_2
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1299__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__253__D tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_tck clkbuf_0_tck/X VGND VGND VPWR VPWR clkbuf_2_3_0_tck/A sky130_fd_sc_hd__clkbuf_1
X__dut__._2714_ clkbuf_5_9_0_tck/X __dut__._2714_/D __dut__._2538_/Y VGND VGND VPWR
+ VPWR __dut__._2714_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2645_ __dut__._2654_/CLK __dut__._2645_/D __dut__._2607_/Y VGND VGND VPWR
+ VPWR __dut__._2645_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2576_ rst VGND VGND VPWR VPWR __dut__._2576_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1527_ _234_/Y __dut__._2688_/Q VGND VGND VPWR VPWR __dut__._1527_/X sky130_fd_sc_hd__and2_4
XFILLER_74_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1458_ __dut__._1466_/A1 __dut__._1456_/X __dut__._1457_/X VGND VGND VPWR
+ VPWR __dut__._2670_/D sky130_fd_sc_hd__a21o_4
XFILLER_34_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1389_ __dut__._2095_/A __dut__._2652_/Q VGND VGND VPWR VPWR __dut__._1389_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2593__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2299__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_268_ _271_/CLK _268_/D VGND VGND VPWR VPWR _268_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_199_ _202_/A VGND VGND VPWR VPWR _199_/X sky130_fd_sc_hd__buf_2
XFILLER_10_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1937__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_162_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1900_ __dut__.__uuf__._1900_/A VGND VGND VPWR VPWR __dut__._2028_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1831_ __dut__.__uuf__._1852_/A __dut__.__uuf__._1831_/B __dut__.__uuf__._1831_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1832_/A sky130_fd_sc_hd__or3_4
XFILLER_33_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1762_ __dut__._1979_/B __dut__._1985_/B __dut__.__uuf__._1761_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1763_/C sky130_fd_sc_hd__o21ai_4
X__dut__.__uuf__._1693_ __dut__._2331_/B __dut__.__uuf__._1688_/X __dut__._2267_/B
+ __dut__.__uuf__._1689_/X VGND VGND VPWR VPWR prod[18] sky130_fd_sc_hd__o22a_4
XFILLER_119_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1847__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1479__A __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2314_ __dut__.__uuf__._2323_/CLK __dut__._2132_/X __dut__.__uuf__._1483_/X
+ VGND VGND VPWR VPWR __dut__._2133_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2245_ __dut__.__uuf__._2288_/CLK __dut__._1994_/X __dut__.__uuf__._1638_/X
+ VGND VGND VPWR VPWR __dut__._1995_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2430_ rst VGND VGND VPWR VPWR __dut__._2430_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2176_ VGND VGND VPWR VPWR __dut__.__uuf__._2176_/HI tie[121] sky130_fd_sc_hd__conb_1
XFILLER_102_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1127_ __dut__.__uuf__._1118_/X __dut__.__uuf__._1114_/X __dut__._2301_/B
+ __dut__._2303_/B __dut__.__uuf__._1126_/X VGND VGND VPWR VPWR __dut__._2300_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_46_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2361_ rst VGND VGND VPWR VPWR __dut__._2361_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1312_ __dut__._1282_/Y mc[16] __dut__._1311_/X VGND VGND VPWR VPWR __dut__._1312_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._2292_ __dut__._2356_/A1 __dut__._2292_/A2 __dut__._2291_/X VGND VGND VPWR
+ VPWR __dut__._2292_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1058_ __dut__.__uuf__._1103_/A VGND VGND VPWR VPWR __dut__.__uuf__._1058_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_28_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1938__A2 prod[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_122_ _312_/Q VGND VGND VPWR VPWR _235_/A sky130_fd_sc_hd__inv_2
XFILLER_137_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1757__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2628_ clkbuf_5_2_0_tck/X __dut__._2628_/D __dut__._2624_/Y VGND VGND VPWR
+ VPWR __dut__._2628_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2588__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2559_ rst VGND VGND VPWR VPWR __dut__._2559_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2314__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_115_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2030_ __dut__._1368_/X VGND VGND VPWR VPWR __dut__.__uuf__._2034_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_111_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2498__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_17_0_tck clkbuf_4_8_0_tck/X VGND VGND VPWR VPWR __dut__._2894_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2290__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1814_ __dut__.__uuf__._1807_/A __dut__.__uuf__._1812_/B __dut__.__uuf__._1782_/X
+ VGND VGND VPWR VPWR __dut__._1994_/A2 sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1745_ __dut__.__uuf__._1768_/A __dut__.__uuf__._1745_/B __dut__.__uuf__._1745_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1746_/A sky130_fd_sc_hd__or3_4
XFILLER_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1930_ __dut__._2328_/A1 prod[22] __dut__._1929_/X VGND VGND VPWR VPWR __dut__._2884_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1577__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1676_ __dut__._2305_/B __dut__.__uuf__._1674_/X __dut__._2241_/B
+ __dut__.__uuf__._1675_/X VGND VGND VPWR VPWR prod[5] sky130_fd_sc_hd__o22a_4
XFILLER_106_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1861_ __dut__._2213_/A __dut__._2849_/Q VGND VGND VPWR VPWR __dut__._1861_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1792_ __dut__._1794_/A1 tie[123] __dut__._1791_/X VGND VGND VPWR VPWR __dut__._2815_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2228_ __dut__.__uuf__._2355_/CLK __dut__._1960_/X __dut__.__uuf__._1658_/X
+ VGND VGND VPWR VPWR __dut__._1961_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_48_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2413_ rst VGND VGND VPWR VPWR __dut__._2413_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2851__CLK clkbuf_5_6_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2159_ VGND VGND VPWR VPWR __dut__.__uuf__._2159_/HI tie[104] sky130_fd_sc_hd__conb_1
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2201__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2344_ __dut__._2356_/A1 __dut__._2344_/A2 __dut__._2343_/X VGND VGND VPWR
+ VPWR __dut__._2344_/X sky130_fd_sc_hd__a21o_4
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_63_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2275_ __dut__._2275_/A __dut__._2275_/B VGND VGND VPWR VPWR __dut__._2275_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_302 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1325_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_313 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1951_/A
+ sky130_fd_sc_hd__buf_2
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_324 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1441_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_335 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2189_/A
+ sky130_fd_sc_hd__buf_2
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1487__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_125_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1530_ __dut__.__uuf__._1522_/X __dut__.__uuf__._1517_/X __dut__._2113_/B
+ __dut__.__uuf__._1527_/X __dut__.__uuf__._1529_/X VGND VGND VPWR VPWR __dut__._2112_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1461_ __dut__.__uuf__._1461_/A VGND VGND VPWR VPWR __dut__.__uuf__._1462_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_143_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1392_ __dut__.__uuf__._1401_/A VGND VGND VPWR VPWR __dut__.__uuf__._1392_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_0_0_tck clkbuf_5_1_0_tck/A VGND VGND VPWR VPWR clkbuf_5_0_0_tck/X sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1838__A1 __dut__._2176_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2013_ __dut__._2071_/B __dut__._2077_/B __dut__.__uuf__._2012_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._2014_/C sky130_fd_sc_hd__o21ai_4
XFILLER_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2060_ __dut__._2060_/A1 __dut__._2060_/A2 __dut__._2059_/X VGND VGND VPWR
+ VPWR __dut__._2060_/X sky130_fd_sc_hd__a21o_4
XFILLER_53_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1728_ __dut__._1328_/X VGND VGND VPWR VPWR __dut__.__uuf__._1732_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_154_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1913_ __dut__._2327_/A __dut__._2875_/Q VGND VGND VPWR VPWR __dut__._1913_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1659_ __dut__.__uuf__._1660_/A VGND VGND VPWR VPWR __dut__.__uuf__._1659_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_146_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2893_ __dut__._2894_/CLK __dut__._2893_/D __dut__._2359_/Y VGND VGND VPWR
+ VPWR __dut__._2893_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1844_ __dut__._1854_/A1 tie[149] __dut__._1843_/X VGND VGND VPWR VPWR __dut__._2841_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_150_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1775_ __dut__._2213_/A __dut__._2806_/Q VGND VGND VPWR VPWR __dut__._1775_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1667__A __dut__._1528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2327_ __dut__._2327_/A __dut__._2327_/B VGND VGND VPWR VPWR __dut__._2327_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2258_ __dut__._2258_/A1 __dut__._2258_/A2 __dut__._2257_/X VGND VGND VPWR
+ VPWR __dut__._2258_/X sky130_fd_sc_hd__a21o_4
XFILLER_140_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_121 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2030_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_110 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1354_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2189_ __dut__._2189_/A __dut__._2189_/B VGND VGND VPWR VPWR __dut__._2189_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_154 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1682_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_132 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1610_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_143 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1624_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_165 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1900_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_176 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2322_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_187 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2356_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_198 psn_inst_psn_buff_203/A VGND VGND VPWR VPWR __dut__._2070_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_129_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1945__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1296__A2 mc[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_242_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1513_ __dut__.__uuf__._1516_/A VGND VGND VPWR VPWR __dut__.__uuf__._1513_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_128_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1444_ __dut__.__uuf__._1270_/X __dut__.__uuf__._1443_/X __dut__._2151_/B
+ __dut__.__uuf__._1270_/X VGND VGND VPWR VPWR __dut__._2150_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1855__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1375_ __dut__.__uuf__._1375_/A VGND VGND VPWR VPWR __dut__.__uuf__._1375_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_89_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1560_ __dut__._1564_/A1 tie[7] __dut__._1559_/X VGND VGND VPWR VPWR __dut__._2699_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1491_ _234_/Y __dut__._2679_/Q VGND VGND VPWR VPWR __dut__._1491_/X sky130_fd_sc_hd__and2_4
XFILLER_100_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2112_ __dut__._2112_/A1 __dut__._2112_/A2 __dut__._2111_/X VGND VGND VPWR
+ VPWR __dut__._2112_/X sky130_fd_sc_hd__a21o_4
XFILLER_14_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2043_ __dut__._2051_/A __dut__._2043_/B VGND VGND VPWR VPWR __dut__._2043_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_26_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_7_0_tck clkbuf_4_7_0_tck/A VGND VGND VPWR VPWR clkbuf_4_7_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2876_ __dut__._2885_/CLK __dut__._2876_/D __dut__._2376_/Y VGND VGND VPWR
+ VPWR __dut__._2876_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1765__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1827_ __dut__._1853_/A __dut__._2832_/Q VGND VGND VPWR VPWR __dut__._1827_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1758_ __dut__._1854_/A1 tie[106] __dut__._1757_/X VGND VGND VPWR VPWR __dut__._2798_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_89_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1689_ __dut__._1689_/A __dut__._2763_/Q VGND VGND VPWR VPWR __dut__._1689_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_3_2_0___dut__.__uuf__.__clk_source___A clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2596__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_192_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1160_ __dut__.__uuf__._1147_/X __dut__.__uuf__._1159_/X __dut__._2279_/B
+ __dut__._2281_/B __dut__.__uuf__._1156_/X VGND VGND VPWR VPWR __dut__._2278_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1091_ __dut__.__uuf__._1149_/A VGND VGND VPWR VPWR __dut__.__uuf__._1102_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_67_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._1993_ __dut__.__uuf__._2014_/A __dut__.__uuf__._1993_/B __dut__.__uuf__._1993_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1994_/A sky130_fd_sc_hd__or3_4
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2730_ __dut__._2744_/CLK __dut__._2730_/D __dut__._2522_/Y VGND VGND VPWR
+ VPWR __dut__._2730_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1585__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2661_ __dut__._2661_/CLK __dut__._2661_/D __dut__._2591_/Y VGND VGND VPWR
+ VPWR __dut__._2661_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1427_ __dut__._2159_/B VGND VGND VPWR VPWR __dut__.__uuf__._1427_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1612_ __dut__._1616_/A1 tie[33] __dut__._1611_/X VGND VGND VPWR VPWR __dut__._2725_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1358_ __dut__.__uuf__._1357_/Y __dut__.__uuf__._1336_/X __dut__.__uuf__._1337_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1358_/X sky130_fd_sc_hd__o21a_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2592_ rst VGND VGND VPWR VPWR __dut__._2592_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1543_ _234_/Y __dut__._2692_/Q VGND VGND VPWR VPWR __dut__._1543_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1289_ __dut__.__uuf__._1281_/Y __dut__.__uuf__._2047_/A __dut__.__uuf__._1283_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1289_/X sky130_fd_sc_hd__o21a_4
XFILLER_105_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1474_ __dut__._1616_/A1 __dut__._1472_/X __dut__._1473_/X VGND VGND VPWR
+ VPWR __dut__._2674_/D sky130_fd_sc_hd__a21o_4
XFILLER_65_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1432__A2 mp[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2026_ __dut__._2030_/A1 __dut__._2026_/A2 __dut__._2025_/X VGND VGND VPWR
+ VPWR __dut__._2026_/X sky130_fd_sc_hd__a21o_4
X_284_ _288_/CLK _284_/D VGND VGND VPWR VPWR _284_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1495__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2859_ clkbuf_5_5_0_tck/X __dut__._2859_/D __dut__._2393_/Y VGND VGND VPWR
+ VPWR __dut__._2859_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_12_0___dut__.__uuf__.__clk_source__ clkbuf_3_6_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2398_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2330_ __dut__.__uuf__._2335_/CLK __dut__._2164_/X __dut__.__uuf__._1407_/X
+ VGND VGND VPWR VPWR __dut__._2165_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2261_ __dut__.__uuf__._2270_/CLK __dut__._2026_/X __dut__.__uuf__._1617_/X
+ VGND VGND VPWR VPWR __dut__._2027_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_114_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1212_ __dut__.__uuf__._1220_/A VGND VGND VPWR VPWR __dut__.__uuf__._1212_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2192_ VGND VGND VPWR VPWR __dut__.__uuf__._2192_/HI tie[137] sky130_fd_sc_hd__conb_1
XFILLER_102_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1143_ __dut__.__uuf__._1146_/A VGND VGND VPWR VPWR __dut__.__uuf__._1143_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_142_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1074_ __dut__.__uuf__._2054_/A VGND VGND VPWR VPWR __dut__.__uuf__._1086_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_28_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1976_ __dut__.__uuf__._1969_/A __dut__.__uuf__._1974_/B __dut__.__uuf__._1944_/X
+ VGND VGND VPWR VPWR __dut__._2054_/A2 sky130_fd_sc_hd__o21a_4
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2808__CLK clkbuf_opt_1_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2713_ __dut__._2721_/CLK __dut__._2713_/D __dut__._2539_/Y VGND VGND VPWR
+ VPWR __dut__._2713_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2644_ __dut__._2654_/CLK __dut__._2644_/D __dut__._2608_/Y VGND VGND VPWR
+ VPWR __dut__._2644_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_psn_inst_psn_buff_93_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2575_ rst VGND VGND VPWR VPWR __dut__._2575_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1526_ __dut__._1530_/A1 __dut__._1524_/X __dut__._1525_/X VGND VGND VPWR
+ VPWR __dut__._2687_/D sky130_fd_sc_hd__a21o_4
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1457_ __dut__._2149_/A __dut__._2669_/Q VGND VGND VPWR VPWR __dut__._1457_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1388_ __dut__._1282_/Y mp[1] __dut__._1387_/X VGND VGND VPWR VPWR __dut__._1388_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_34_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._2009_ __dut__._2213_/A __dut__._2009_/B VGND VGND VPWR VPWR __dut__._2009_/X
+ sky130_fd_sc_hd__and2_4
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_267_ _271_/CLK _267_/D VGND VGND VPWR VPWR _267_/Q sky130_fd_sc_hd__dfxtp_4
X_198_ _198_/A VGND VGND VPWR VPWR _198_/X sky130_fd_sc_hd__buf_2
XFILLER_115_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1892__A2 prod[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_155_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2243__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_322_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1830_ __dut__._2003_/B __dut__._2009_/B __dut__.__uuf__._1829_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1831_/C sky130_fd_sc_hd__o21ai_4
XFILLER_33_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1761_ __dut__.__uuf__._1761_/A VGND VGND VPWR VPWR __dut__.__uuf__._1761_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1692_ __dut__._2329_/B __dut__.__uuf__._1688_/X __dut__._2265_/B
+ __dut__.__uuf__._1689_/X VGND VGND VPWR VPWR prod[17] sky130_fd_sc_hd__o22a_4
XFILLER_146_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2313_ __dut__.__uuf__._2323_/CLK __dut__._2130_/X __dut__.__uuf__._1488_/X
+ VGND VGND VPWR VPWR __dut__._2131_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2244_ __dut__.__uuf__._2282_/CLK __dut__._1992_/X __dut__.__uuf__._1639_/X
+ VGND VGND VPWR VPWR __dut__._1993_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1863__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1332__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2175_ VGND VGND VPWR VPWR __dut__.__uuf__._2175_/HI tie[120] sky130_fd_sc_hd__conb_1
XFILLER_102_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1495__A __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1126_ __dut__.__uuf__._1141_/A VGND VGND VPWR VPWR __dut__.__uuf__._1126_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2360_ rst VGND VGND VPWR VPWR __dut__._2360_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1311_ _234_/Y __dut__._2634_/Q VGND VGND VPWR VPWR __dut__._1311_/X sky130_fd_sc_hd__and2_4
X__dut__._2291_ __dut__._2313_/A __dut__._2291_/B VGND VGND VPWR VPWR __dut__._2291_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1057_ __dut__.__uuf__._1057_/A VGND VGND VPWR VPWR __dut__.__uuf__._1057_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_83_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1959_ __dut__._2051_/B __dut__._2057_/B __dut__.__uuf__._1958_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1960_/C sky130_fd_sc_hd__o21ai_4
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_121_ _289_/Q VGND VGND VPWR VPWR _230_/A sky130_fd_sc_hd__buf_2
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1773__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2627_ clkbuf_5_3_0_tck/X __dut__._2627_/D __dut__._2625_/Y VGND VGND VPWR
+ VPWR __dut__._2627_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2558_ rst VGND VGND VPWR VPWR __dut__._2558_/Y sky130_fd_sc_hd__inv_2
X__dut__._1509_ __dut__._1617_/A __dut__._2681_/Q VGND VGND VPWR VPWR __dut__._1509_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2489_ rst VGND VGND VPWR VPWR __dut__._2489_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_272_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_tck clkbuf_0_tck/X VGND VGND VPWR VPWR clkbuf_2_1_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_61_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1813_ __dut__.__uuf__._1813_/A VGND VGND VPWR VPWR __dut__._1996_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_139_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1744_ __dut__.__uuf__._1276_/X __dut__.__uuf__._1742_/B __dut__.__uuf__._1742_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1745_/C sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1675_ __dut__.__uuf__._1682_/A VGND VGND VPWR VPWR __dut__.__uuf__._1675_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_146_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1860_ __dut__._1860_/A1 tie[157] __dut__._1859_/X VGND VGND VPWR VPWR __dut__._2849_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1791_ __dut__._1793_/A __dut__._2814_/Q VGND VGND VPWR VPWR __dut__._1791_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2289__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1593__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2227_ __dut__.__uuf__._2355_/CLK __dut__._1958_/X __dut__.__uuf__._1659_/X
+ VGND VGND VPWR VPWR __dut__._1959_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_130_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2412_ rst VGND VGND VPWR VPWR __dut__._2412_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2158_ VGND VGND VPWR VPWR __dut__.__uuf__._2158_/HI tie[103] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2089_ VGND VGND VPWR VPWR __dut__.__uuf__._2089_/HI tie[34] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1109_ __dut__.__uuf__._1103_/X __dut__.__uuf__._1100_/X __dut__._2313_/B
+ __dut__._2315_/B __dut__.__uuf__._1097_/X VGND VGND VPWR VPWR __dut__._2312_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._2343_ __dut__._2349_/A __dut__._2343_/B VGND VGND VPWR VPWR __dut__._2343_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_29_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2274_ __dut__._2274_/A1 __dut__._2274_/A2 __dut__._2273_/X VGND VGND VPWR
+ VPWR __dut__._2274_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_56_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_303 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1313_/A
+ sky130_fd_sc_hd__buf_2
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_314 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1549_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_325 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2149_/A
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_336 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2227_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_24_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1544__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1989_ __dut__._2213_/A __dut__._1989_/B VGND VGND VPWR VPWR __dut__._1989_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_112_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2599__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2024__A __dut__.__uuf__._2044_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_118_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1460_ __dut__.__uuf__._1472_/A VGND VGND VPWR VPWR __dut__.__uuf__._1460_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1391_ __dut__.__uuf__._1378_/X __dut__.__uuf__._1390_/X __dut__._2173_/B
+ __dut__.__uuf__._1378_/X VGND VGND VPWR VPWR __dut__._2172_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2012_ __dut__.__uuf__._2012_/A VGND VGND VPWR VPWR __dut__.__uuf__._2012_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1727_ __dut__._1963_/B __dut__.__uuf__._1725_/X __dut__._1962_/A2
+ VGND VGND VPWR VPWR __dut__._1964_/A2 sky130_fd_sc_hd__a21boi_4
XFILLER_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1912_ __dut__._2328_/A1 prod[13] __dut__._1911_/X VGND VGND VPWR VPWR __dut__._2875_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2892_ __dut__._2892_/CLK __dut__._2892_/D __dut__._2360_/Y VGND VGND VPWR
+ VPWR __dut__._2892_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1658_ __dut__.__uuf__._1660_/A VGND VGND VPWR VPWR __dut__.__uuf__._1658_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1843_ __dut__._1853_/A __dut__._2840_/Q VGND VGND VPWR VPWR __dut__._1843_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2699__CLK clkbuf_5_2_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1589_ __dut__.__uuf__._1593_/A VGND VGND VPWR VPWR __dut__.__uuf__._1589_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1774_ __dut__._1774_/A1 tie[114] __dut__._1773_/X VGND VGND VPWR VPWR __dut__._2806_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2326_ __dut__._2328_/A1 __dut__._2326_/A2 __dut__._2325_/X VGND VGND VPWR
+ VPWR __dut__._2326_/X sky130_fd_sc_hd__a21o_4
X__dut__._2257_ __dut__._2257_/A __dut__._2257_/B VGND VGND VPWR VPWR __dut__._2257_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2304__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_111 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1358_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_100 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2108_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2188_ __dut__._2200_/A1 __dut__._2188_/A2 __dut__._2187_/X VGND VGND VPWR
+ VPWR __dut__._2188_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_144 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1626_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_133 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1602_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_155 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1684_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_122 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1952_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_166 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1722_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_188 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2328_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_177 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2266_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_129_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_16_0_tck clkbuf_4_8_0_tck/X VGND VGND VPWR VPWR __dut__._2744_/CLK sky130_fd_sc_hd__clkbuf_1
Xpsn_inst_psn_buff_199 psn_inst_psn_buff_203/A VGND VGND VPWR VPWR __dut__._2064_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_144_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1961__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_235_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__265__CLK _270_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1756__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2841__CLK clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1512_ __dut__.__uuf__._1501_/X __dut__.__uuf__._1495_/X __dut__._2121_/B
+ __dut__.__uuf__._1506_/X __dut__.__uuf__._1511_/X VGND VGND VPWR VPWR __dut__._2120_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1508__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1443_ __dut__.__uuf__._1442_/Y __dut__.__uuf__._1438_/X __dut__.__uuf__._1337_/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._1443_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1374_ __dut__.__uuf__._1367_/X __dut__.__uuf__._1373_/X __dut__._2179_/B
+ __dut__.__uuf__._1367_/X VGND VGND VPWR VPWR __dut__._2178_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1871__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1490_ __dut__._1490_/A1 __dut__._1488_/X __dut__._1489_/X VGND VGND VPWR
+ VPWR __dut__._2678_/D sky130_fd_sc_hd__a21o_4
XFILLER_100_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2111_ __dut__._2111_/A __dut__._2111_/B VGND VGND VPWR VPWR __dut__._2111_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2042_ __dut__._2044_/A1 __dut__._2042_/A2 __dut__._2041_/X VGND VGND VPWR
+ VPWR __dut__._2042_/X sky130_fd_sc_hd__a21o_4
XFILLER_110_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2207__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_19_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2875_ __dut__._2885_/CLK __dut__._2875_/D __dut__._2377_/Y VGND VGND VPWR
+ VPWR __dut__._2875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1826_ __dut__._1854_/A1 tie[140] __dut__._1825_/X VGND VGND VPWR VPWR __dut__._2832_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2172__A1 __dut__._2176_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1757_ __dut__._1853_/A __dut__._2797_/Q VGND VGND VPWR VPWR __dut__._1757_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1781__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1688_ __dut__._1688_/A1 tie[71] __dut__._1687_/X VGND VGND VPWR VPWR __dut__._2763_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_95_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2309_ __dut__._2313_/A __dut__._2309_/B VGND VGND VPWR VPWR __dut__._2309_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_44_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2117__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_185_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1090_ __dut__.__uuf__._1655_/A VGND VGND VPWR VPWR __dut__.__uuf__._1149_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1992_ __dut__._2063_/B __dut__._2069_/B __dut__.__uuf__._1991_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1993_/C sky130_fd_sc_hd__o21ai_4
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2660_ clkbuf_5_3_0_tck/X __dut__._2660_/D __dut__._2592_/Y VGND VGND VPWR
+ VPWR __dut__._2660_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1498__A __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1426_ __dut__.__uuf__._1426_/A VGND VGND VPWR VPWR __dut__.__uuf__._1426_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1611_ __dut__._1611_/A __dut__._2724_/Q VGND VGND VPWR VPWR __dut__._1611_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1357_ __dut__._2187_/B VGND VGND VPWR VPWR __dut__.__uuf__._1357_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._2591_ rst VGND VGND VPWR VPWR __dut__._2591_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1542_ __dut__._1542_/A1 __dut__._1540_/X __dut__._1541_/X VGND VGND VPWR
+ VPWR __dut__._2691_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1288_ __dut__.__uuf__._1507_/A VGND VGND VPWR VPWR __dut__.__uuf__._2047_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_46_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1473_ __dut__._1473_/A __dut__._2673_/Q VGND VGND VPWR VPWR __dut__._1473_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_105_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2025_ __dut__._2029_/A __dut__._2025_/B VGND VGND VPWR VPWR __dut__._2025_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_139_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_283_ _288_/CLK _283_/D VGND VGND VPWR VPWR _283_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2858_ clkbuf_5_4_0_tck/X __dut__._2858_/D __dut__._2394_/Y VGND VGND VPWR
+ VPWR __dut__._2858_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1809_ __dut__._2213_/A __dut__._2823_/Q VGND VGND VPWR VPWR __dut__._1809_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2789_ _308_/CLK __dut__._2789_/D __dut__._2463_/Y VGND VGND VPWR VPWR __dut__._2789_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_150_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2400__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_100_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_9_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_145_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2260_ __dut__.__uuf__._2270_/CLK __dut__._2024_/X __dut__.__uuf__._1620_/X
+ VGND VGND VPWR VPWR __dut__._2025_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_141_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1211_ __dut__.__uuf__._1207_/X __dut__.__uuf__._1204_/X __dut__._2245_/B
+ __dut__._2247_/B __dut__.__uuf__._1200_/X VGND VGND VPWR VPWR __dut__._2244_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._2191_ VGND VGND VPWR VPWR __dut__.__uuf__._2191_/HI tie[136] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1142_ __dut__.__uuf__._1133_/X __dut__.__uuf__._1130_/X __dut__._2291_/B
+ __dut__._2293_/B __dut__.__uuf__._1141_/X VGND VGND VPWR VPWR __dut__._2290_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_28_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1073_ __dut__.__uuf__._1072_/X __dut__.__uuf__._1069_/X __dut__._2337_/B
+ __dut__._2339_/B __dut__.__uuf__._1066_/X VGND VGND VPWR VPWR __dut__._2336_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_83_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_6_0_tck clkbuf_4_7_0_tck/A VGND VGND VPWR VPWR clkbuf_4_6_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1975_ __dut__.__uuf__._1975_/A VGND VGND VPWR VPWR __dut__._2056_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2712_ __dut__._2721_/CLK __dut__._2712_/D __dut__._2540_/Y VGND VGND VPWR
+ VPWR __dut__._2712_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1409_ __dut__.__uuf__._1408_/Y __dut__.__uuf__._1388_/X __dut__.__uuf__._1389_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1409_/X sky130_fd_sc_hd__o21a_4
XFILLER_78_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2643_ __dut__._2661_/CLK __dut__._2643_/D __dut__._2609_/Y VGND VGND VPWR
+ VPWR __dut__._2643_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2389_ __dut__.__uuf__._2426_/CLK __dut__._2282_/X __dut__.__uuf__._1152_/X
+ VGND VGND VPWR VPWR __dut__._2283_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_132_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2574_ rst VGND VGND VPWR VPWR __dut__._2574_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1525_ __dut__._1525_/A __dut__._2686_/Q VGND VGND VPWR VPWR __dut__._1525_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_86_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1456_ __dut__._1282_/Y mp[17] __dut__._1455_/X VGND VGND VPWR VPWR __dut__._1456_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_92_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1387_ _234_/Y __dut__._2653_/Q VGND VGND VPWR VPWR __dut__._1387_/X sky130_fd_sc_hd__and2_4
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2008_ __dut__._2008_/A1 __dut__._2008_/A2 __dut__._2007_/X VGND VGND VPWR
+ VPWR __dut__._2008_/X sky130_fd_sc_hd__a21o_4
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_266_ _270_/CLK _266_/D VGND VGND VPWR VPWR _266_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_197_ _198_/A VGND VGND VPWR VPWR _197_/X sky130_fd_sc_hd__buf_2
XFILLER_142_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_148_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_315_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1760_ __dut__._1979_/B __dut__._1985_/B VGND VGND VPWR VPWR __dut__.__uuf__._1761_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1691_ __dut__._2327_/B __dut__.__uuf__._1688_/X __dut__._2263_/B
+ __dut__.__uuf__._1689_/X VGND VGND VPWR VPWR prod[16] sky130_fd_sc_hd__o22a_4
XFILLER_20_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2305__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2312_ __dut__.__uuf__._2323_/CLK __dut__._2128_/X __dut__.__uuf__._1491_/X
+ VGND VGND VPWR VPWR __dut__._2129_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_88_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2243_ __dut__.__uuf__._2282_/CLK __dut__._1990_/X __dut__.__uuf__._1640_/X
+ VGND VGND VPWR VPWR __dut__._1991_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_153_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1332__A2 mc[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2174_ VGND VGND VPWR VPWR __dut__.__uuf__._2174_/HI tie[119] sky130_fd_sc_hd__conb_1
XFILLER_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1125_ __dut__.__uuf__._1132_/A VGND VGND VPWR VPWR __dut__.__uuf__._1125_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_68_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1310_ __dut__._1346_/A1 __dut__._1308_/X __dut__._1309_/X VGND VGND VPWR
+ VPWR __dut__._2633_/D sky130_fd_sc_hd__a21o_4
XFILLER_110_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2290_ __dut__._2356_/A1 __dut__._2290_/A2 __dut__._2289_/X VGND VGND VPWR
+ VPWR __dut__._2290_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1056_ __dut__.__uuf__._1034_/X __dut__.__uuf__._1055_/X __dut__._2349_/B
+ __dut__._2351_/B __dut__.__uuf__._1051_/X VGND VGND VPWR VPWR __dut__._2348_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_83_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__291__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1958_ __dut__.__uuf__._1958_/A VGND VGND VPWR VPWR __dut__.__uuf__._1958_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_120_ _308_/Q VGND VGND VPWR VPWR _120_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1889_ __dut__.__uuf__._1889_/A VGND VGND VPWR VPWR __dut__._2024_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2348__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2626_ rst VGND VGND VPWR VPWR __dut__._2626_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2557_ rst VGND VGND VPWR VPWR __dut__._2557_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__308__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1508_ __dut__._1282_/Y mp[28] __dut__._1507_/X VGND VGND VPWR VPWR __dut__._1508_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._2488_ rst VGND VGND VPWR VPWR __dut__._2488_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1439_ _234_/Y __dut__._2666_/Q VGND VGND VPWR VPWR __dut__._1439_/X sky130_fd_sc_hd__and2_4
XFILLER_61_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_249_ _197_/X _249_/D VGND VGND VPWR VPWR _249_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_143_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2125__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_265_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2360__CLK __dut__.__uuf__._2402_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1812_ __dut__.__uuf__._1823_/A __dut__.__uuf__._1812_/B __dut__.__uuf__._1812_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1813_/A sky130_fd_sc_hd__or3_4
XFILLER_40_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1743_ __dut__.__uuf__._1743_/A VGND VGND VPWR VPWR __dut__.__uuf__._1745_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_147_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1674_ __dut__.__uuf__._1681_/A VGND VGND VPWR VPWR __dut__.__uuf__._1674_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_20_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1790_ __dut__._1790_/A1 tie[122] __dut__._1789_/X VGND VGND VPWR VPWR __dut__._2814_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2226_ __dut__.__uuf__._2355_/CLK __dut__._1956_/X __dut__.__uuf__._1660_/X
+ VGND VGND VPWR VPWR __dut__._1957_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2411_ rst VGND VGND VPWR VPWR __dut__._2411_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2157_ VGND VGND VPWR VPWR __dut__.__uuf__._2157_/HI tie[102] sky130_fd_sc_hd__conb_1
XFILLER_57_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2088_ VGND VGND VPWR VPWR __dut__.__uuf__._2088_/HI tie[33] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1108_ __dut__.__uuf__._1116_/A VGND VGND VPWR VPWR __dut__.__uuf__._1108_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2342_ __dut__._2342_/A1 __dut__._2342_/A2 __dut__._2341_/X VGND VGND VPWR
+ VPWR __dut__._2342_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1039_ __dut__.__uuf__._1191_/A VGND VGND VPWR VPWR __dut__.__uuf__._1244_/A
+ sky130_fd_sc_hd__inv_2
X__dut__._2273_ __dut__._2273_/A __dut__._2273_/B VGND VGND VPWR VPWR __dut__._2273_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_113_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_304 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1309_/A
+ sky130_fd_sc_hd__buf_2
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_315 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1793_/A
+ sky130_fd_sc_hd__buf_8
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_337 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2239_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_326 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1953_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA_psn_inst_psn_buff_49_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2233__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1544__A2 mc[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1988_ __dut__._2000_/A1 __dut__._1988_/A2 __dut__._1987_/X VGND VGND VPWR
+ VPWR __dut__._1988_/X sky130_fd_sc_hd__a21o_4
XFILLER_152_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2609_ rst VGND VGND VPWR VPWR __dut__._2609_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1480__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1959__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1390_ __dut__.__uuf__._1387_/Y __dut__.__uuf__._1388_/X __dut__.__uuf__._1389_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1390_/X sky130_fd_sc_hd__o21a_4
XFILLER_143_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2011_ __dut__._2071_/B __dut__._2077_/B VGND VGND VPWR VPWR __dut__.__uuf__._2012_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_69_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1869__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1726_ __dut__._1963_/B __dut__.__uuf__._1725_/X __dut__.__uuf__._1998_/A
+ VGND VGND VPWR VPWR __dut__._1962_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1911_ __dut__._2327_/A __dut__._2874_/Q VGND VGND VPWR VPWR __dut__._1911_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_5_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2891_ __dut__._2892_/CLK __dut__._2891_/D __dut__._2361_/Y VGND VGND VPWR
+ VPWR __dut__._2891_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1657_ __dut__.__uuf__._1660_/A VGND VGND VPWR VPWR __dut__.__uuf__._1657_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1842_ __dut__._2176_/A1 tie[148] __dut__._1841_/X VGND VGND VPWR VPWR __dut__._2840_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1588_ __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR __dut__.__uuf__._1593_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1773_ __dut__._2213_/A __dut__._2805_/Q VGND VGND VPWR VPWR __dut__._1773_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_150_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2209_ VGND VGND VPWR VPWR __dut__.__uuf__._2209_/HI tie[154] sky130_fd_sc_hd__conb_1
XFILLER_124_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2325_ __dut__._2325_/A __dut__._2325_/B VGND VGND VPWR VPWR __dut__._2325_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2256_ __dut__._2256_/A1 __dut__._2256_/A2 __dut__._2255_/X VGND VGND VPWR
+ VPWR __dut__._2256_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_112 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1346_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_101 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2106_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._2187_ __dut__._2189_/A __dut__._2187_/B VGND VGND VPWR VPWR __dut__._2187_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1779__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_134 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1790_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_145 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1644_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_123 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1548_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_167 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1902_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_189 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2256_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_156 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1694_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_178 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2268_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1204__A __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2403__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2793__CLK _270_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1961__B __dut__._1961_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_130_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2279__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_148_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1511_ __dut__._1456_/X __dut__.__uuf__._1502_/X __dut__._2123_/B
+ __dut__.__uuf__._1507_/X VGND VGND VPWR VPWR __dut__.__uuf__._1511_/X sky130_fd_sc_hd__o22a_4
XFILLER_156_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1508__A2 mp[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1442_ __dut__._2153_/B VGND VGND VPWR VPWR __dut__.__uuf__._1442_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_143_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1373_ __dut__.__uuf__._1372_/Y __dut__.__uuf__._1362_/X __dut__.__uuf__._1363_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1373_/X sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._2313__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1784__A __dut__._1532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2110_ __dut__._2110_/A1 __dut__._2110_/A2 __dut__._2109_/X VGND VGND VPWR
+ VPWR __dut__._2110_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1444__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2041_ __dut__._2051_/A __dut__._2041_/B VGND VGND VPWR VPWR __dut__._2041_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_110_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1599__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1709_ __dut__._2355_/B __dut__.__uuf__._1681_/A __dut__._2291_/B
+ __dut__.__uuf__._1682_/A VGND VGND VPWR VPWR prod[30] sky130_fd_sc_hd__o22a_4
XFILLER_126_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2874_ __dut__._2885_/CLK __dut__._2874_/D __dut__._2378_/Y VGND VGND VPWR
+ VPWR __dut__._2874_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1825_ __dut__._1853_/A __dut__._2831_/Q VGND VGND VPWR VPWR __dut__._1825_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1756_ __dut__._1854_/A1 tie[105] __dut__._1755_/X VGND VGND VPWR VPWR __dut__._2797_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_135_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1687_ __dut__._1687_/A __dut__._2762_/Q VGND VGND VPWR VPWR __dut__._1687_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_2_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2308_ __dut__._2356_/A1 __dut__._2308_/A2 __dut__._2307_/X VGND VGND VPWR
+ VPWR __dut__._2308_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2239_ __dut__._2239_/A __dut__._2239_/B VGND VGND VPWR VPWR __dut__._2239_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_32_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2133__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_178_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1674__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1991_ __dut__.__uuf__._1991_/A VGND VGND VPWR VPWR __dut__.__uuf__._1991_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_63_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2689__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1425_ __dut__.__uuf__._1418_/X __dut__.__uuf__._1424_/X __dut__._2159_/B
+ __dut__.__uuf__._1418_/X VGND VGND VPWR VPWR __dut__._2158_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1610_ __dut__._1610_/A1 tie[32] __dut__._1609_/X VGND VGND VPWR VPWR __dut__._2724_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1356_ __dut__.__uuf__._1375_/A VGND VGND VPWR VPWR __dut__.__uuf__._1356_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2590_ rst VGND VGND VPWR VPWR __dut__._2590_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1541_ __dut__._1541_/A __dut__._2690_/Q VGND VGND VPWR VPWR __dut__._1541_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1287_ __dut__.__uuf__._1307_/A VGND VGND VPWR VPWR __dut__.__uuf__._1507_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_86_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1472_ __dut__._1282_/Y mp[20] __dut__._1471_/X VGND VGND VPWR VPWR __dut__._1472_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_105_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_15_0_tck clkbuf_4_7_0_tck/X VGND VGND VPWR VPWR __dut__._2680_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_42_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2024_ __dut__._2024_/A1 __dut__._2024_/A2 __dut__._2023_/X VGND VGND VPWR
+ VPWR __dut__._2024_/X sky130_fd_sc_hd__a21o_4
XFILLER_139_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_282_ _288_/CLK _282_/D VGND VGND VPWR VPWR _282_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_31_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1689__A __dut__._1528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2857_ clkbuf_5_4_0_tck/X __dut__._2857_/D __dut__._2395_/Y VGND VGND VPWR
+ VPWR __dut__._2857_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1808_ __dut__._1810_/A1 tie[131] __dut__._1807_/X VGND VGND VPWR VPWR __dut__._2823_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2788_ __dut__._2885_/CLK __dut__._2788_/D __dut__._2464_/Y VGND VGND VPWR
+ VPWR __dut__._2788_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1739_ __dut__._2327_/A __dut__._2788_/Q VGND VGND VPWR VPWR __dut__._1739_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA__255__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2831__CLK __dut__._2845_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1408__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1967__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2317__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_145_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_295_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1210_ __dut__.__uuf__._1220_/A VGND VGND VPWR VPWR __dut__.__uuf__._1210_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2190_ VGND VGND VPWR VPWR __dut__.__uuf__._2190_/HI tie[135] sky130_fd_sc_hd__conb_1
XFILLER_141_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1141_ __dut__.__uuf__._1141_/A VGND VGND VPWR VPWR __dut__.__uuf__._1141_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1072_ __dut__.__uuf__._1103_/A VGND VGND VPWR VPWR __dut__.__uuf__._1072_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1974_ __dut__.__uuf__._1985_/A __dut__.__uuf__._1974_/B __dut__.__uuf__._1974_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1975_/A sky130_fd_sc_hd__or3_4
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1877__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2711_ clkbuf_5_8_0_tck/X __dut__._2711_/D __dut__._2541_/Y VGND VGND VPWR
+ VPWR __dut__._2711_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1408_ __dut__._2167_/B VGND VGND VPWR VPWR __dut__.__uuf__._1408_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_116_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2642_ __dut__._2661_/CLK __dut__._2642_/D __dut__._2610_/Y VGND VGND VPWR
+ VPWR __dut__._2642_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1886__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2388_ __dut__.__uuf__._2415_/CLK __dut__._2280_/X __dut__.__uuf__._1154_/X
+ VGND VGND VPWR VPWR __dut__._2281_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2854__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1339_ __dut__.__uuf__._1326_/X __dut__.__uuf__._1338_/X __dut__._2193_/B
+ __dut__.__uuf__._1326_/X VGND VGND VPWR VPWR __dut__._2192_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._2573_ rst VGND VGND VPWR VPWR __dut__._2573_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2501__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1524_ __dut__._1282_/Y start __dut__._1523_/X VGND VGND VPWR VPWR __dut__._1524_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_79_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1455_ _234_/Y __dut__._2670_/Q VGND VGND VPWR VPWR __dut__._1455_/X sky130_fd_sc_hd__and2_4
XFILLER_27_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1386_ __dut__._1386_/A1 __dut__._1384_/X __dut__._1385_/X VGND VGND VPWR
+ VPWR __dut__._2652_/D sky130_fd_sc_hd__a21o_4
XFILLER_92_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2007_ __dut__._2213_/A __dut__._2007_/B VGND VGND VPWR VPWR __dut__._2007_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_265_ _270_/CLK _265_/D VGND VGND VPWR VPWR _265_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1787__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_196_ _198_/A VGND VGND VPWR VPWR _196_/X sky130_fd_sc_hd__buf_2
XFILLER_41_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2411__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_210_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_308_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1690_ __dut__._2325_/B __dut__.__uuf__._1688_/X __dut__._2261_/B
+ __dut__.__uuf__._1689_/X VGND VGND VPWR VPWR prod[15] sky130_fd_sc_hd__o22a_4
XFILLER_118_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2311_ __dut__.__uuf__._2323_/CLK __dut__._2126_/X __dut__.__uuf__._1494_/X
+ VGND VGND VPWR VPWR __dut__._2127_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2242_ __dut__.__uuf__._2282_/CLK __dut__._1988_/X __dut__.__uuf__._1641_/X
+ VGND VGND VPWR VPWR __dut__._1989_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2173_ VGND VGND VPWR VPWR __dut__.__uuf__._2173_/HI tie[118] sky130_fd_sc_hd__conb_1
XFILLER_99_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1124_ __dut__.__uuf__._1118_/X __dut__.__uuf__._1114_/X __dut__._2303_/B
+ __dut__._2305_/B __dut__.__uuf__._1111_/X VGND VGND VPWR VPWR __dut__._2302_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1055_ __dut__.__uuf__._1114_/A VGND VGND VPWR VPWR __dut__.__uuf__._1055_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1957_ __dut__._2051_/B __dut__._2057_/B VGND VGND VPWR VPWR __dut__.__uuf__._1958_/A
+ sky130_fd_sc_hd__and2_4
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1888_ __dut__.__uuf__._1931_/A __dut__.__uuf__._1888_/B __dut__.__uuf__._1888_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1889_/A sky130_fd_sc_hd__or3_4
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2231__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2625_ rst VGND VGND VPWR VPWR __dut__._2625_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2556_ rst VGND VGND VPWR VPWR __dut__._2556_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2487_ rst VGND VGND VPWR VPWR __dut__._2487_/Y sky130_fd_sc_hd__inv_2
X__dut__._1507_ _234_/Y __dut__._2683_/Q VGND VGND VPWR VPWR __dut__._1507_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2284__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1438_ __dut__._1442_/A1 __dut__._1436_/X __dut__._1437_/X VGND VGND VPWR
+ VPWR __dut__._2665_/D sky130_fd_sc_hd__a21o_4
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1369_ __dut__._2095_/A __dut__._2647_/Q VGND VGND VPWR VPWR __dut__._1369_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1207__A __dut__.__uuf__._1478_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2406__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_248_ _198_/X _312_/Q VGND VGND VPWR VPWR _248_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_179_ _270_/Q _186_/B VGND VGND VPWR VPWR _269_/D sky130_fd_sc_hd__or2_4
XFILLER_143_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_tck clkbuf_4_5_0_tck/A VGND VGND VPWR VPWR clkbuf_4_5_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2141__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_160_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_258_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1811_ __dut__.__uuf__._1766_/X __dut__.__uuf__._1809_/B __dut__.__uuf__._1809_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1812_/C sky130_fd_sc_hd__o21a_4
XFILLER_61_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1742_ __dut__.__uuf__._1742_/A __dut__.__uuf__._1742_/B __dut__.__uuf__._1742_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1743_/A sky130_fd_sc_hd__or3_4
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1673_ __dut__._2303_/B __dut__.__uuf__._1666_/X __dut__._2239_/B
+ __dut__.__uuf__._1668_/X VGND VGND VPWR VPWR prod[4] sky130_fd_sc_hd__o22a_4
XFILLER_146_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2225_ __dut__.__uuf__._2402_/CLK __dut__._1954_/X __dut__.__uuf__._1661_/X
+ VGND VGND VPWR VPWR __dut__._1955_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2410_ rst VGND VGND VPWR VPWR __dut__._2410_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2156_ VGND VGND VPWR VPWR __dut__.__uuf__._2156_/HI tie[101] sky130_fd_sc_hd__conb_1
XFILLER_57_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1107_ __dut__.__uuf__._1103_/X __dut__.__uuf__._1100_/X __dut__._2315_/B
+ __dut__._2317_/B __dut__.__uuf__._1097_/X VGND VGND VPWR VPWR __dut__._2314_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_113_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2087_ VGND VGND VPWR VPWR __dut__.__uuf__._2087_/HI tie[32] sky130_fd_sc_hd__conb_1
X__dut__._2341_ __dut__._2341_/A __dut__._2341_/B VGND VGND VPWR VPWR __dut__._2341_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2272_ __dut__._2272_/A1 __dut__._2272_/A2 __dut__._2271_/X VGND VGND VPWR
+ VPWR __dut__._2272_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1038_ __dut__.__uuf__._1998_/A VGND VGND VPWR VPWR __dut__.__uuf__._1038_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_113_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_316 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1611_/A
+ sky130_fd_sc_hd__buf_4
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_338 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1701_/A
+ sky130_fd_sc_hd__buf_2
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_305 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1305_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_327 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2221_/A
+ sky130_fd_sc_hd__buf_2
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1987_ __dut__._2213_/A __dut__._1987_/B VGND VGND VPWR VPWR __dut__._1987_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2608_ rst VGND VGND VPWR VPWR __dut__._2608_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2539_ rst VGND VGND VPWR VPWR __dut__._2539_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1480__A2 mp[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1975__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2010_ __dut__._1360_/X VGND VGND VPWR VPWR __dut__.__uuf__._2014_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_112_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1725_ __dut__._2215_/B __dut__._1380_/X VGND VGND VPWR VPWR __dut__.__uuf__._1725_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_119_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1910_ __dut__._1910_/A1 prod[12] __dut__._1909_/X VGND VGND VPWR VPWR __dut__._2874_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2890_ __dut__._2892_/CLK __dut__._2890_/D __dut__._2362_/Y VGND VGND VPWR
+ VPWR __dut__._2890_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1656_ __dut__.__uuf__._1660_/A VGND VGND VPWR VPWR __dut__.__uuf__._1656_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1841_ __dut__._2213_/A __dut__._2839_/Q VGND VGND VPWR VPWR __dut__._1841_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1885__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1587_ __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR __dut__.__uuf__._1612_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_108_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1772_ __dut__._1772_/A1 tie[113] __dut__._1771_/X VGND VGND VPWR VPWR __dut__._2805_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_103_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2208_ VGND VGND VPWR VPWR __dut__.__uuf__._2208_/HI tie[153] sky130_fd_sc_hd__conb_1
XFILLER_102_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2139_ VGND VGND VPWR VPWR __dut__.__uuf__._2139_/HI tie[84] sky130_fd_sc_hd__conb_1
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2324_ __dut__._2324_/A1 __dut__._2324_/A2 __dut__._2323_/X VGND VGND VPWR
+ VPWR __dut__._2324_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_61_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2255_ __dut__._2255_/A __dut__._2255_/B VGND VGND VPWR VPWR __dut__._2255_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_102 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2104_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._2186_ __dut__._2200_/A1 __dut__._2186_/A2 __dut__._2185_/X VGND VGND VPWR
+ VPWR __dut__._2186_/X sky130_fd_sc_hd__a21o_4
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_135 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1554_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_146 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1646_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_124 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1578_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_113 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1322_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_168 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1904_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_157 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1690_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_179 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2270_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_40_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1795__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2350__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_98_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__.__uuf__._1890__A __dut__.__uuf__._1890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_123_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1510_ __dut__.__uuf__._1516_/A VGND VGND VPWR VPWR __dut__.__uuf__._1510_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1441_ __dut__.__uuf__._1449_/A VGND VGND VPWR VPWR __dut__.__uuf__._1441_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1372_ __dut__._2181_/B VGND VGND VPWR VPWR __dut__.__uuf__._1372_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_143_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1444__A2 mp[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2040_ __dut__._2046_/A1 __dut__._2040_/A2 __dut__._2039_/X VGND VGND VPWR
+ VPWR __dut__._2040_/X sky130_fd_sc_hd__a21o_4
XFILLER_110_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1708_ __dut__._2353_/B __dut__.__uuf__._1702_/X __dut__._2289_/B
+ __dut__.__uuf__._1703_/X VGND VGND VPWR VPWR prod[29] sky130_fd_sc_hd__o22a_4
XFILLER_119_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1639_ __dut__.__uuf__._1642_/A VGND VGND VPWR VPWR __dut__.__uuf__._1639_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2504__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2873_ __dut__._2885_/CLK __dut__._2873_/D __dut__._2379_/Y VGND VGND VPWR
+ VPWR __dut__._2873_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1824_ __dut__._1854_/A1 tie[139] __dut__._1823_/X VGND VGND VPWR VPWR __dut__._2831_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_123_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1040__A __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1755_ __dut__._1853_/A __dut__._2796_/Q VGND VGND VPWR VPWR __dut__._1755_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1380__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1686_ __dut__._1688_/A1 tie[70] __dut__._1685_/X VGND VGND VPWR VPWR __dut__._2762_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2307_ __dut__._2313_/A __dut__._2307_/B VGND VGND VPWR VPWR __dut__._2307_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2238_ __dut__._2238_/A1 __dut__._2238_/A2 __dut__._2237_/X VGND VGND VPWR
+ VPWR __dut__._2238_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1215__A __dut__.__uuf__._1215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2169_ __dut__._2189_/A __dut__._2169_/B VGND VGND VPWR VPWR __dut__._2169_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2414__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_240_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_338_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2246__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_82_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1990_ __dut__._2063_/B __dut__._2069_/B VGND VGND VPWR VPWR __dut__.__uuf__._1991_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1424_ __dut__.__uuf__._1423_/Y __dut__.__uuf__._1413_/X __dut__.__uuf__._1414_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1424_/X sky130_fd_sc_hd__o21a_4
XFILLER_144_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1355_ __dut__.__uuf__._1355_/A VGND VGND VPWR VPWR __dut__.__uuf__._1375_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_132_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1540_ __dut__._1282_/Y mc[8] __dut__._1539_/X VGND VGND VPWR VPWR __dut__._1540_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1286_ __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR __dut__.__uuf__._1286_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1471_ _234_/Y __dut__._2674_/Q VGND VGND VPWR VPWR __dut__._1471_/X sky130_fd_sc_hd__and2_4
XFILLER_73_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1403__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2023_ __dut__._2029_/A __dut__._2023_/B VGND VGND VPWR VPWR __dut__._2023_/X
+ sky130_fd_sc_hd__and2_4
X_281_ _288_/CLK _281_/D VGND VGND VPWR VPWR _281_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_psn_inst_psn_buff_24_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2856_ clkbuf_5_5_0_tck/X __dut__._2856_/D __dut__._2396_/Y VGND VGND VPWR
+ VPWR __dut__._2856_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1807_ __dut__._2213_/A __dut__._2822_/Q VGND VGND VPWR VPWR __dut__._1807_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2787_ __dut__._2892_/CLK __dut__._2787_/D __dut__._2465_/Y VGND VGND VPWR
+ VPWR __dut__._2787_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1738_ __dut__._2328_/A1 tie[96] __dut__._1737_/X VGND VGND VPWR VPWR __dut__._2788_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1669_ __dut__._1673_/A __dut__._2753_/Q VGND VGND VPWR VPWR __dut__._1669_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_18_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1408__A2 mp[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2409__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_190_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_288_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1983__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1344__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1140_ __dut__.__uuf__._1146_/A VGND VGND VPWR VPWR __dut__.__uuf__._1140_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1071_ __dut__.__uuf__._1071_/A VGND VGND VPWR VPWR __dut__.__uuf__._1071_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1973_ __dut__.__uuf__._1929_/X __dut__.__uuf__._1971_/B __dut__.__uuf__._1971_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1974_/C sky130_fd_sc_hd__o21a_4
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2710_ clkbuf_5_8_0_tck/X __dut__._2710_/D __dut__._2542_/Y VGND VGND VPWR
+ VPWR __dut__._2710_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2641_ __dut__._2357_/B __dut__._2641_/D __dut__._2611_/Y VGND VGND VPWR
+ VPWR __dut__._2641_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1407_ __dut__.__uuf__._1426_/A VGND VGND VPWR VPWR __dut__.__uuf__._1407_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_116_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1886__A2 prod[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2387_ __dut__.__uuf__._2415_/CLK __dut__._2278_/X __dut__.__uuf__._1158_/X
+ VGND VGND VPWR VPWR __dut__._2279_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_104_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1338_ __dut__.__uuf__._1334_/Y __dut__.__uuf__._1336_/X __dut__.__uuf__._1337_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1338_/X sky130_fd_sc_hd__o21a_4
X__dut__._2572_ rst VGND VGND VPWR VPWR __dut__._2572_/Y sky130_fd_sc_hd__inv_2
X__dut__._1523_ _234_/Y __dut__._2687_/Q VGND VGND VPWR VPWR __dut__._1523_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1269_ __dut__.__uuf__._1269_/A VGND VGND VPWR VPWR __dut__.__uuf__._1269_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1454_ __dut__._1454_/A1 __dut__._1452_/X __dut__._1453_/X VGND VGND VPWR
+ VPWR __dut__._2669_/D sky130_fd_sc_hd__a21o_4
XFILLER_92_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1385_ __dut__._2095_/A __dut__._2651_/Q VGND VGND VPWR VPWR __dut__._1385_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2229__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2006_ __dut__._2008_/A1 __dut__._2006_/A2 __dut__._2005_/X VGND VGND VPWR
+ VPWR __dut__._2006_/X sky130_fd_sc_hd__a21o_4
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_264_ _270_/CLK _264_/D VGND VGND VPWR VPWR _264_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_195_ _198_/A VGND VGND VPWR VPWR _195_/X sky130_fd_sc_hd__buf_2
XFILLER_127_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2839_ clkbuf_opt_2_tck/A __dut__._2839_/D __dut__._2413_/Y VGND VGND VPWR
+ VPWR __dut__._2839_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2139__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_14_0_tck clkbuf_4_7_0_tck/X VGND VGND VPWR VPWR __dut__._2726_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2310_ __dut__.__uuf__._2323_/CLK __dut__._2124_/X __dut__.__uuf__._1500_/X
+ VGND VGND VPWR VPWR __dut__._2125_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_127_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2241_ __dut__.__uuf__._2282_/CLK __dut__._1986_/X __dut__.__uuf__._1642_/X
+ VGND VGND VPWR VPWR __dut__._1987_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_142_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2602__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2172_ VGND VGND VPWR VPWR __dut__.__uuf__._2172_/HI tie[117] sky130_fd_sc_hd__conb_1
Xclkbuf_5_29_0_tck clkbuf_5_29_0_tck/A VGND VGND VPWR VPWR clkbuf_opt_2_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_101_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1123_ __dut__.__uuf__._1132_/A VGND VGND VPWR VPWR __dut__.__uuf__._1123_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1054_ __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR __dut__.__uuf__._1114_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1956_ __dut__._1340_/X VGND VGND VPWR VPWR __dut__.__uuf__._1960_/B
+ sky130_fd_sc_hd__inv_2
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_1_1_0_tck_A clkbuf_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1887_ __dut__.__uuf__._1875_/X __dut__.__uuf__._1885_/B __dut__.__uuf__._1885_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1888_/C sky130_fd_sc_hd__o21a_4
XFILLER_137_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1308__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2512__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2624_ rst VGND VGND VPWR VPWR __dut__._2624_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2555_ rst VGND VGND VPWR VPWR __dut__._2555_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_91_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1506_ __dut__._1506_/A1 __dut__._1504_/X __dut__._1505_/X VGND VGND VPWR
+ VPWR __dut__._2682_/D sky130_fd_sc_hd__a21o_4
XFILLER_143_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2486_ rst VGND VGND VPWR VPWR __dut__._2486_/Y sky130_fd_sc_hd__inv_2
X__dut__._1437_ __dut__._1441_/A __dut__._2664_/Q VGND VGND VPWR VPWR __dut__._1437_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2307__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1368_ __dut__._1282_/Y mc[29] __dut__._1367_/X VGND VGND VPWR VPWR __dut__._1368_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1299_ _234_/Y __dut__._2631_/Q VGND VGND VPWR VPWR __dut__._1299_/X sky130_fd_sc_hd__and2_4
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_247_ _199_/X _311_/Q VGND VGND VPWR VPWR _247_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__.__uuf__._1223__A __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_178_ _271_/Q _181_/B VGND VGND VPWR VPWR _270_/D sky130_fd_sc_hd__and2_4
XFILLER_143_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2422__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2054__A __dut__.__uuf__._2054_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_153_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_320_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1810_ __dut__.__uuf__._1810_/A VGND VGND VPWR VPWR __dut__.__uuf__._1812_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA__268__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1741_ __dut__._1971_/B __dut__._1977_/B __dut__.__uuf__._1740_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1742_/C sky130_fd_sc_hd__o21ai_4
XANTENNA___dut__._2844__CLK __dut__._2845_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1672_ __dut__._2301_/B __dut__.__uuf__._1666_/X __dut__._2237_/B
+ __dut__.__uuf__._1668_/X VGND VGND VPWR VPWR prod[3] sky130_fd_sc_hd__o22a_4
XANTENNA___dut__.__uuf__._1133__A __dut__.__uuf__._1177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2224_ VGND VGND VPWR VPWR __dut__.__uuf__._2224_/HI tie[169] sky130_fd_sc_hd__conb_1
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2155_ VGND VGND VPWR VPWR __dut__.__uuf__._2155_/HI tie[100] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._1710__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1106_ __dut__.__uuf__._1116_/A VGND VGND VPWR VPWR __dut__.__uuf__._1106_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_113_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2086_ VGND VGND VPWR VPWR __dut__.__uuf__._2086_/HI tie[31] sky130_fd_sc_hd__conb_1
X__dut__._2340_ __dut__._2340_/A1 __dut__._2340_/A2 __dut__._2339_/X VGND VGND VPWR
+ VPWR __dut__._2340_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1037_ __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR __dut__.__uuf__._1998_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._2271_ __dut__._2271_/A __dut__._2271_/B VGND VGND VPWR VPWR __dut__._2271_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpsn_inst_psn_buff_317 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1555_/A
+ sky130_fd_sc_hd__buf_2
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_306 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1301_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_328 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2219_/A
+ sky130_fd_sc_hd__buf_2
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2507__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_339 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2251_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1939_ __dut__.__uuf__._1960_/A __dut__.__uuf__._1939_/B __dut__.__uuf__._1939_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1940_/A sky130_fd_sc_hd__or3_4
XFILLER_24_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1411__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1986_ __dut__._2000_/A1 __dut__._1986_/A2 __dut__._1985_/X VGND VGND VPWR
+ VPWR __dut__._1986_/X sky130_fd_sc_hd__a21o_4
XFILLER_140_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2607_ rst VGND VGND VPWR VPWR __dut__._2607_/Y sky130_fd_sc_hd__inv_2
X__dut__._2538_ rst VGND VGND VPWR VPWR __dut__._2538_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2469_ rst VGND VGND VPWR VPWR __dut__._2469_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1218__A __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2417__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_270_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1991__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2327__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1724_ __dut__.__uuf__._1716_/A __dut__.__uuf__._1721_/B __dut__.__uuf__._1723_/X
+ VGND VGND VPWR VPWR __dut__._1958_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_119_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1655_ __dut__.__uuf__._1655_/A VGND VGND VPWR VPWR __dut__.__uuf__._1660_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1840_ __dut__._2176_/A1 tie[147] __dut__._1839_/X VGND VGND VPWR VPWR __dut__._2839_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_147_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1586_ __dut__.__uuf__._1586_/A VGND VGND VPWR VPWR __dut__.__uuf__._1586_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1771_ __dut__._2213_/A __dut__._2804_/Q VGND VGND VPWR VPWR __dut__._1771_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_108_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2207_ VGND VGND VPWR VPWR __dut__.__uuf__._2207_/HI tie[152] sky130_fd_sc_hd__conb_1
XFILLER_0_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2138_ VGND VGND VPWR VPWR __dut__.__uuf__._2138_/HI tie[83] sky130_fd_sc_hd__conb_1
XFILLER_75_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2069_ VGND VGND VPWR VPWR __dut__.__uuf__._2069_/HI tie[14] sky130_fd_sc_hd__conb_1
X__dut__._2323_ __dut__._2323_/A __dut__._2323_/B VGND VGND VPWR VPWR __dut__._2323_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1038__A __dut__.__uuf__._1998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2254_ __dut__._2256_/A1 __dut__._2254_/A2 __dut__._2253_/X VGND VGND VPWR
+ VPWR __dut__._2254_/X sky130_fd_sc_hd__a21o_4
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_103 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2102_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._2185_ __dut__._2189_/A __dut__._2185_/B VGND VGND VPWR VPWR __dut__._2185_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_54_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_125 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1580_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_114 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1318_/A1
+ sky130_fd_sc_hd__buf_2
Xclkbuf_4_4_0_tck clkbuf_4_5_0_tck/A VGND VGND VPWR VPWR clkbuf_5_9_0_tck/A sky130_fd_sc_hd__clkbuf_1
Xpsn_inst_psn_buff_136 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2036_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_147 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1660_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_169 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1906_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_158 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1688_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_149_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1501__A __dut__.__uuf__._1564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1969_ __dut__._2213_/A __dut__._1969_/B VGND VGND VPWR VPWR __dut__._1969_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2051__B __dut__._1957_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_116_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1440_ __dut__.__uuf__._1429_/X __dut__.__uuf__._1439_/X __dut__._2153_/B
+ __dut__.__uuf__._1429_/X VGND VGND VPWR VPWR __dut__._2152_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1371_ __dut__.__uuf__._1375_/A VGND VGND VPWR VPWR __dut__.__uuf__._1371_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_104_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_0_0_tck_A clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2610__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0___dut__.__uuf__.__clk_source__ clkbuf_4_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2348_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2057__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1707_ __dut__._2351_/B __dut__.__uuf__._1702_/X __dut__._2287_/B
+ __dut__.__uuf__._1703_/X VGND VGND VPWR VPWR prod[28] sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1638_ __dut__.__uuf__._1642_/A VGND VGND VPWR VPWR __dut__.__uuf__._1638_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2872_ __dut__._2885_/CLK __dut__._2872_/D __dut__._2380_/Y VGND VGND VPWR
+ VPWR __dut__._2872_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1823_ __dut__._1853_/A __dut__._2830_/Q VGND VGND VPWR VPWR __dut__._1823_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_119_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1569_ __dut__._1396_/X __dut__.__uuf__._1565_/X __dut__._2095_/B
+ __dut__.__uuf__._1309_/A VGND VGND VPWR VPWR __dut__.__uuf__._1569_/X sky130_fd_sc_hd__o22a_4
XFILLER_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1754_ __dut__._1854_/A1 tie[104] __dut__._1753_/X VGND VGND VPWR VPWR __dut__._2796_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1380__A2 mc[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2520__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1685_ __dut__._1685_/A __dut__._2761_/Q VGND VGND VPWR VPWR __dut__._1685_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_135_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2306_ __dut__._2356_/A1 __dut__._2306_/A2 __dut__._2305_/X VGND VGND VPWR
+ VPWR __dut__._2306_/X sky130_fd_sc_hd__a21o_4
XFILLER_29_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2237_ __dut__._2239_/A __dut__._2237_/B VGND VGND VPWR VPWR __dut__._2237_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2168_ __dut__._2180_/A1 __dut__._2168_/A2 __dut__._2167_/X VGND VGND VPWR
+ VPWR __dut__._2168_/X sky130_fd_sc_hd__a21o_4
X__dut__._2099_ __dut__._2099_/A __dut__._2099_/B VGND VGND VPWR VPWR __dut__._2099_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2430__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_233_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2605__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1423_ __dut__._2161_/B VGND VGND VPWR VPWR __dut__.__uuf__._1423_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_144_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1354_ __dut__.__uuf__._1342_/X __dut__.__uuf__._1352_/X __dut__._2187_/B
+ __dut__.__uuf__._1353_/X VGND VGND VPWR VPWR __dut__._2186_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1285_ __dut__.__uuf__._1295_/A VGND VGND VPWR VPWR __dut__.__uuf__._1285_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_98_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1470_ __dut__._1616_/A1 __dut__._1468_/X __dut__._1469_/X VGND VGND VPWR
+ VPWR __dut__._2673_/D sky130_fd_sc_hd__a21o_4
XFILLER_86_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2022_ __dut__._2024_/A1 __dut__._2022_/A2 __dut__._2021_/X VGND VGND VPWR
+ VPWR __dut__._2022_/X sky130_fd_sc_hd__a21o_4
XFILLER_42_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_280_ _288_/CLK _280_/D VGND VGND VPWR VPWR _280_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__.__uuf__._1035__B __dut__._1957_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_17_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2515__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1051__A __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2855_ clkbuf_5_5_0_tck/X __dut__._2855_/D __dut__._2397_/Y VGND VGND VPWR
+ VPWR __dut__._2855_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1806_ __dut__._1806_/A1 tie[130] __dut__._1805_/X VGND VGND VPWR VPWR __dut__._2822_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2786_ __dut__._2885_/CLK __dut__._2786_/D __dut__._2466_/Y VGND VGND VPWR
+ VPWR __dut__._2786_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1737_ __dut__._2327_/A __dut__._2787_/Q VGND VGND VPWR VPWR __dut__._1737_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2302__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1668_ __dut__._1668_/A1 tie[61] __dut__._1667_/X VGND VGND VPWR VPWR __dut__._2753_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_92_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1599_ __dut__._1793_/A __dut__._2718_/Q VGND VGND VPWR VPWR __dut__._1599_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_91_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2425__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1344__A2 mc[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_183_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1070_ __dut__.__uuf__._1058_/X __dut__.__uuf__._1069_/X __dut__._2339_/B
+ __dut__._2341_/B __dut__.__uuf__._1066_/X VGND VGND VPWR VPWR __dut__._2338_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_95_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2363__CLK __dut__.__uuf__._2402_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1972_ __dut__.__uuf__._1972_/A VGND VGND VPWR VPWR __dut__.__uuf__._1974_/B
+ sky130_fd_sc_hd__inv_2
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2640_ __dut__._2357_/B __dut__._2640_/D __dut__._2612_/Y VGND VGND VPWR
+ VPWR __dut__._2640_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2386_ __dut__.__uuf__._2415_/CLK __dut__._2276_/X __dut__.__uuf__._1161_/X
+ VGND VGND VPWR VPWR __dut__._2277_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1406_ __dut__.__uuf__._1476_/A VGND VGND VPWR VPWR __dut__.__uuf__._1426_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_120_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1337_ __dut__.__uuf__._1337_/A VGND VGND VPWR VPWR __dut__.__uuf__._1337_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_116_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2571_ rst VGND VGND VPWR VPWR __dut__._2571_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1522_ __dut__._1530_/A1 __dut__._1520_/X __dut__._1521_/X VGND VGND VPWR
+ VPWR __dut__._2686_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1268_ __dut__.__uuf__._1263_/B __dut__.__uuf__._1266_/X __dut__.__uuf__._1229_/X
+ __dut__._2219_/B __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR __dut__._2218_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_74_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1453_ __dut__._2149_/A __dut__._2668_/Q VGND VGND VPWR VPWR __dut__._1453_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1199_ __dut__.__uuf__._1206_/A VGND VGND VPWR VPWR __dut__.__uuf__._1199_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1384_ __dut__._1282_/Y mp[0] __dut__._1383_/X VGND VGND VPWR VPWR __dut__._1384_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_54_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2005_ __dut__._2213_/A __dut__._2005_/B VGND VGND VPWR VPWR __dut__._2005_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_42_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_263_ _193_/A _263_/D VGND VGND VPWR VPWR _263_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_194_ _202_/A VGND VGND VPWR VPWR _198_/A sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2236__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2838_ clkbuf_opt_2_tck/X __dut__._2838_/D __dut__._2414_/Y VGND VGND VPWR
+ VPWR __dut__._2838_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2769_ __dut__._2865_/CLK __dut__._2769_/D __dut__._2483_/Y VGND VGND VPWR
+ VPWR __dut__._2769_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2240_ __dut__.__uuf__._2282_/CLK __dut__._1984_/X __dut__.__uuf__._1644_/X
+ VGND VGND VPWR VPWR __dut__._1985_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2171_ VGND VGND VPWR VPWR __dut__.__uuf__._2171_/HI tie[116] sky130_fd_sc_hd__conb_1
XFILLER_102_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1122_ __dut__.__uuf__._1118_/X __dut__.__uuf__._1114_/X __dut__._2305_/B
+ __dut__._2307_/B __dut__.__uuf__._1111_/X VGND VGND VPWR VPWR __dut__._2304_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1053_ __dut__.__uuf__._1057_/A VGND VGND VPWR VPWR __dut__.__uuf__._1053_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_56_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1955_ __dut__.__uuf__._1948_/A __dut__.__uuf__._1953_/B __dut__.__uuf__._1944_/X
+ VGND VGND VPWR VPWR __dut__._2046_/A2 sky130_fd_sc_hd__o21a_4
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1886_ __dut__.__uuf__._1886_/A VGND VGND VPWR VPWR __dut__.__uuf__._1888_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_137_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2065__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1308__A2 mc[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2623_ rst VGND VGND VPWR VPWR __dut__._2623_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2369_ __dut__.__uuf__._2372_/CLK __dut__._2242_/X __dut__.__uuf__._1212_/X
+ VGND VGND VPWR VPWR __dut__._2243_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_120_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2554_ rst VGND VGND VPWR VPWR __dut__._2554_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1505_ __dut__._1505_/A __dut__._2671_/Q VGND VGND VPWR VPWR __dut__._1505_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_84_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2485_ rst VGND VGND VPWR VPWR __dut__._2485_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1436_ __dut__._1282_/Y mp[12] __dut__._1435_/X VGND VGND VPWR VPWR __dut__._1436_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1492__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1367_ _234_/Y __dut__._2648_/Q VGND VGND VPWR VPWR __dut__._1367_/X sky130_fd_sc_hd__and2_4
X__dut__._1298_ __dut__._1564_/A1 __dut__._1296_/X __dut__._1297_/X VGND VGND VPWR
+ VPWR __dut__._2630_/D sky130_fd_sc_hd__a21o_4
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_246_ _200_/X _310_/Q VGND VGND VPWR VPWR _246_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_177_ _272_/Q _181_/B VGND VGND VPWR VPWR _271_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2796__CLK _270_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1319__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_146_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1989__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_313_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2401__CLK __dut__.__uuf__._2402_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1740_ __dut__.__uuf__._1740_/A VGND VGND VPWR VPWR __dut__.__uuf__._1740_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_119_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1671_ __dut__._2299_/B __dut__.__uuf__._1666_/X __dut__._2235_/B
+ __dut__.__uuf__._1668_/X VGND VGND VPWR VPWR prod[2] sky130_fd_sc_hd__o22a_4
Xclkbuf_3_0_0___dut__.__uuf__.__clk_source__ clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_1_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_107_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2613__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2223_ VGND VGND VPWR VPWR __dut__.__uuf__._2223_/HI tie[168] sky130_fd_sc_hd__conb_1
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2154_ VGND VGND VPWR VPWR __dut__.__uuf__._2154_/HI tie[99] sky130_fd_sc_hd__conb_1
XFILLER_130_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1105_ __dut__.__uuf__._1149_/A VGND VGND VPWR VPWR __dut__.__uuf__._1116_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2085_ VGND VGND VPWR VPWR __dut__.__uuf__._2085_/HI tie[30] sky130_fd_sc_hd__conb_1
XFILLER_113_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1036_ __dut__.__uuf__._1456_/A VGND VGND VPWR VPWR __dut__.__uuf__._1479_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._2270_ __dut__._2270_/A1 __dut__._2270_/A2 __dut__._2269_/X VGND VGND VPWR
+ VPWR __dut__._2270_/X sky130_fd_sc_hd__a21o_4
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_307 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1297_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_318 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2029_/A
+ sky130_fd_sc_hd__buf_4
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1938_ __dut__._2043_/B __dut__._2049_/B __dut__.__uuf__._1937_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1939_/C sky130_fd_sc_hd__o21ai_4
Xpsn_inst_psn_buff_329 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2217_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_156_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1869_ __dut__._1304_/X VGND VGND VPWR VPWR __dut__.__uuf__._1873_/B
+ sky130_fd_sc_hd__inv_2
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1985_ __dut__._2213_/A __dut__._1985_/B VGND VGND VPWR VPWR __dut__._1985_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2523__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2606_ rst VGND VGND VPWR VPWR __dut__._2606_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2537_ rst VGND VGND VPWR VPWR __dut__._2537_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2468_ rst VGND VGND VPWR VPWR __dut__._2468_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1419_ _234_/Y __dut__._2661_/Q VGND VGND VPWR VPWR __dut__._1419_/X sky130_fd_sc_hd__and2_4
Xclkbuf_5_13_0_tck clkbuf_4_6_0_tck/X VGND VGND VPWR VPWR __dut__._2654_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__._2399_ rst VGND VGND VPWR VPWR __dut__._2399_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_5_28_0_tck clkbuf_5_29_0_tck/A VGND VGND VPWR VPWR _271_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_229_ _229_/A _302_/Q VGND VGND VPWR VPWR _301_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1052__A2 __dut__.__uuf__._1038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2433__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1940__A2 prod[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_263_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1456__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2608__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1723_ __dut__.__uuf__._1890_/A VGND VGND VPWR VPWR __dut__.__uuf__._1723_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_138_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1654_ __dut__.__uuf__._1654_/A VGND VGND VPWR VPWR __dut__.__uuf__._1654_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_119_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1585_ __dut__.__uuf__._1586_/A VGND VGND VPWR VPWR __dut__.__uuf__._1585_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1770_ __dut__._1770_/A1 tie[112] __dut__._1769_/X VGND VGND VPWR VPWR __dut__._2804_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2206_ VGND VGND VPWR VPWR __dut__.__uuf__._2206_/HI tie[151] sky130_fd_sc_hd__conb_1
XFILLER_103_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2137_ VGND VGND VPWR VPWR __dut__.__uuf__._2137_/HI tie[82] sky130_fd_sc_hd__conb_1
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2068_ VGND VGND VPWR VPWR __dut__.__uuf__._2068_/HI tie[13] sky130_fd_sc_hd__conb_1
X__dut__._2322_ __dut__._2322_/A1 __dut__._2322_/A2 __dut__._2321_/X VGND VGND VPWR
+ VPWR __dut__._2322_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2253_ __dut__._2255_/A __dut__._2253_/B VGND VGND VPWR VPWR __dut__._2253_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2518__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2184_ __dut__._2184_/A1 __dut__._2184_/A2 __dut__._2183_/X VGND VGND VPWR
+ VPWR __dut__._2184_/X sky130_fd_sc_hd__a21o_4
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_126 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1584_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_137 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2118_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_104 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2100_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_115 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1506_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA_psn_inst_psn_buff_47_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_148 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1662_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_159 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._2238_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1054__A __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1968_ __dut__._2078_/A1 __dut__._1968_/A2 __dut__._1967_/X VGND VGND VPWR
+ VPWR __dut__._1968_/X sky130_fd_sc_hd__a21o_4
XFILLER_140_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1899_ __dut__._1899_/A __dut__._2868_/Q VGND VGND VPWR VPWR __dut__._1899_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2834__CLK __dut__._2845_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1229__A __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2428__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_109_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__301__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1370_ __dut__.__uuf__._1367_/X __dut__.__uuf__._1369_/X __dut__._2181_/B
+ __dut__.__uuf__._1367_/X VGND VGND VPWR VPWR __dut__._2180_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1507__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2707__CLK clkbuf_5_0_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1706_ __dut__._2349_/B __dut__.__uuf__._1702_/X __dut__._2285_/B
+ __dut__.__uuf__._1703_/X VGND VGND VPWR VPWR prod[27] sky130_fd_sc_hd__o22a_4
XFILLER_135_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2871_ __dut__._2885_/CLK __dut__._2871_/D __dut__._2381_/Y VGND VGND VPWR
+ VPWR __dut__._2871_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1637_ __dut__.__uuf__._1643_/A VGND VGND VPWR VPWR __dut__.__uuf__._1642_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2073__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1822_ __dut__._1854_/A1 tie[138] __dut__._1821_/X VGND VGND VPWR VPWR __dut__._2830_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_119_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1568_ __dut__.__uuf__._1577_/A VGND VGND VPWR VPWR __dut__.__uuf__._1568_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2857__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1753_ __dut__._1853_/A __dut__._2795_/Q VGND VGND VPWR VPWR __dut__._1753_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1499_ __dut__.__uuf__._1581_/A VGND VGND VPWR VPWR __dut__.__uuf__._1516_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_122_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1684_ __dut__._1684_/A1 tie[69] __dut__._1683_/X VGND VGND VPWR VPWR __dut__._2761_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_135_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2305_ __dut__._2313_/A __dut__._2305_/B VGND VGND VPWR VPWR __dut__._2305_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1840__A1 __dut__._2176_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2893__D __dut__._2893_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2236_ __dut__._2238_/A1 __dut__._2236_/A2 __dut__._2235_/X VGND VGND VPWR
+ VPWR __dut__._2236_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2167_ __dut__._2167_/A __dut__._2167_/B VGND VGND VPWR VPWR __dut__._2167_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2098_ __dut__._2098_/A1 __dut__._2098_/A2 __dut__._2097_/X VGND VGND VPWR
+ VPWR __dut__._2098_/X sky130_fd_sc_hd__a21o_4
XFILLER_138_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1327__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1997__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2292__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1422_ __dut__.__uuf__._1426_/A VGND VGND VPWR VPWR __dut__.__uuf__._1422_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_116_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2621__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1353_ __dut__.__uuf__._1393_/A VGND VGND VPWR VPWR __dut__.__uuf__._1353_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_3_0_tck clkbuf_4_3_0_tck/A VGND VGND VPWR VPWR clkbuf_5_7_0_tck/A sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1284_ __dut__.__uuf__._1281_/Y __dut__.__uuf__._2050_/B __dut__.__uuf__._1283_/X
+ VGND VGND VPWR VPWR __dut__._2212_/A2 sky130_fd_sc_hd__o21ai_4
XFILLER_100_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1822__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__294__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2021_ __dut__._2029_/A __dut__._2021_/B VGND VGND VPWR VPWR __dut__._2021_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2854_ clkbuf_5_4_0_tck/X __dut__._2854_/D __dut__._2398_/Y VGND VGND VPWR
+ VPWR __dut__._2854_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1805_ __dut__._2213_/A __dut__._2821_/Q VGND VGND VPWR VPWR __dut__._1805_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2785_ __dut__._2885_/CLK __dut__._2785_/D __dut__._2467_/Y VGND VGND VPWR
+ VPWR __dut__._2785_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2531__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1736_ __dut__._2328_/A1 tie[95] __dut__._1735_/X VGND VGND VPWR VPWR __dut__._2787_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1667_ __dut__._1667_/A __dut__._2752_/Q VGND VGND VPWR VPWR __dut__._1667_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1598_ __dut__._1790_/A1 tie[26] __dut__._1597_/X VGND VGND VPWR VPWR __dut__._2718_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2219_ __dut__._2219_/A __dut__._2219_/B VGND VGND VPWR VPWR __dut__._2219_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_60_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__126__A tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2441__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_176_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1971_ __dut__.__uuf__._2014_/A __dut__.__uuf__._1971_/B __dut__.__uuf__._1971_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1972_/A sky130_fd_sc_hd__or3_4
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2616__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2385_ __dut__.__uuf__._2422_/CLK __dut__._2274_/X __dut__.__uuf__._1166_/X
+ VGND VGND VPWR VPWR __dut__._2275_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1405_ __dut__.__uuf__._1393_/X __dut__.__uuf__._1403_/X __dut__._2167_/B
+ __dut__.__uuf__._1404_/X VGND VGND VPWR VPWR __dut__._2166_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1336_ __dut__.__uuf__._1711_/A VGND VGND VPWR VPWR __dut__.__uuf__._1336_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_120_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2570_ rst VGND VGND VPWR VPWR __dut__._2570_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1521_ __dut__._1521_/A __dut__._2685_/Q VGND VGND VPWR VPWR __dut__._1521_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1267_ __dut__.__uuf__._1341_/A VGND VGND VPWR VPWR __dut__.__uuf__._1326_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2296__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1452_ __dut__._1282_/Y mp[16] __dut__._1451_/X VGND VGND VPWR VPWR __dut__._1452_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1198_ __dut__.__uuf__._1192_/X __dut__.__uuf__._1188_/X __dut__._2253_/B
+ __dut__._2255_/B __dut__.__uuf__._1185_/X VGND VGND VPWR VPWR __dut__._2252_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1383_ _234_/Y __dut__._2652_/Q VGND VGND VPWR VPWR __dut__._1383_/X sky130_fd_sc_hd__and2_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2526__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2004_ __dut__._2008_/A1 __dut__._2004_/A2 __dut__._2003_/X VGND VGND VPWR
+ VPWR __dut__._2004_/X sky130_fd_sc_hd__a21o_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_262_ _193_/A _262_/D VGND VGND VPWR VPWR _262_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_193_ _193_/A VGND VGND VPWR VPWR _202_/A sky130_fd_sc_hd__inv_2
XFILLER_10_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2837_ __dut__._2845_/CLK __dut__._2837_/D __dut__._2415_/Y VGND VGND VPWR
+ VPWR __dut__._2837_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2768_ __dut__._2865_/CLK __dut__._2768_/D __dut__._2484_/Y VGND VGND VPWR
+ VPWR __dut__._2768_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1719_ __dut__._1729_/A __dut__._2778_/Q VGND VGND VPWR VPWR __dut__._1719_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2699_ clkbuf_5_2_0_tck/X __dut__._2699_/D __dut__._2553_/Y VGND VGND VPWR
+ VPWR __dut__._2699_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1605__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2436__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_293_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2170_ VGND VGND VPWR VPWR __dut__.__uuf__._2170_/HI tie[115] sky130_fd_sc_hd__conb_1
XFILLER_114_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1121_ __dut__.__uuf__._1132_/A VGND VGND VPWR VPWR __dut__.__uuf__._1121_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_68_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2278__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1052_ __dut__.__uuf__._1034_/X __dut__.__uuf__._1038_/X __dut__._2351_/B
+ __dut__._2353_/B __dut__.__uuf__._1051_/X VGND VGND VPWR VPWR __dut__._2350_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1515__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1147__A __dut__.__uuf__._1177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1954_ __dut__.__uuf__._1954_/A VGND VGND VPWR VPWR __dut__._2048_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_51_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1885_ __dut__.__uuf__._1906_/A __dut__.__uuf__._1885_/B __dut__.__uuf__._1885_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1886_/A sky130_fd_sc_hd__or3_4
XFILLER_137_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2081__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2622_ rst VGND VGND VPWR VPWR __dut__._2622_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2368_ __dut__.__uuf__._2372_/CLK __dut__._2240_/X __dut__.__uuf__._1214_/X
+ VGND VGND VPWR VPWR __dut__._2241_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1319_ __dut__.__uuf__._1323_/A VGND VGND VPWR VPWR __dut__.__uuf__._1319_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2553_ rst VGND VGND VPWR VPWR __dut__._2553_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2299_ __dut__.__uuf__._2319_/CLK __dut__._2102_/X __dut__.__uuf__._1547_/X
+ VGND VGND VPWR VPWR __dut__._2103_/B sky130_fd_sc_hd__dfrtp_4
Xclkbuf_opt_2_tck clkbuf_opt_2_tck/A VGND VGND VPWR VPWR clkbuf_opt_2_tck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_47_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1504_ __dut__._1282_/Y mc[5] __dut__._1503_/X VGND VGND VPWR VPWR __dut__._1504_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_101_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2484_ rst VGND VGND VPWR VPWR __dut__._2484_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_77_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1492__A2 mp[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1435_ _234_/Y __dut__._2665_/Q VGND VGND VPWR VPWR __dut__._1435_/X sky130_fd_sc_hd__and2_4
XFILLER_15_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1366_ __dut__._1366_/A1 __dut__._1364_/X __dut__._1365_/X VGND VGND VPWR
+ VPWR __dut__._2647_/D sky130_fd_sc_hd__a21o_4
XFILLER_34_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1297_ __dut__._1297_/A __dut__._2629_/Q VGND VGND VPWR VPWR __dut__._1297_/X
+ sky130_fd_sc_hd__and2_4
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_245_ _201_/X _309_/Q VGND VGND VPWR VPWR _245_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_176_ _273_/Q _181_/B VGND VGND VPWR VPWR _272_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2353__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_115_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1335__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_139_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_306_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1670_ __dut__._2297_/B __dut__.__uuf__._1666_/X __dut__._2233_/B
+ __dut__.__uuf__._1668_/X VGND VGND VPWR VPWR prod[1] sky130_fd_sc_hd__o22a_4
XFILLER_146_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2222_ VGND VGND VPWR VPWR __dut__.__uuf__._2222_/HI tie[167] sky130_fd_sc_hd__conb_1
XFILLER_114_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2153_ VGND VGND VPWR VPWR __dut__.__uuf__._2153_/HI tie[98] sky130_fd_sc_hd__conb_1
XFILLER_87_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1104_ __dut__.__uuf__._1103_/X __dut__.__uuf__._1100_/X __dut__._2317_/B
+ __dut__._2319_/B __dut__.__uuf__._1097_/X VGND VGND VPWR VPWR __dut__._2316_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2084_ VGND VGND VPWR VPWR __dut__.__uuf__._2084_/HI tie[29] sky130_fd_sc_hd__conb_1
XFILLER_113_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1035_ __dut__._1955_/B __dut__._1957_/B VGND VGND VPWR VPWR __dut__.__uuf__._1456_/A
+ sky130_fd_sc_hd__or2_4
XANTENNA___dut__.__uuf__._2226__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_319 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1541_/A
+ sky130_fd_sc_hd__buf_2
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_308 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1563_/A
+ sky130_fd_sc_hd__buf_2
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1937_ __dut__.__uuf__._1937_/A VGND VGND VPWR VPWR __dut__.__uuf__._1937_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_138_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1868_ __dut__.__uuf__._1861_/A __dut__.__uuf__._1866_/B __dut__.__uuf__._1836_/X
+ VGND VGND VPWR VPWR __dut__._2014_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_149_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1799_ __dut__.__uuf__._1799_/A VGND VGND VPWR VPWR __dut__.__uuf__._1801_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._1984_ __dut__._2000_/A1 __dut__._1984_/A2 __dut__._1983_/X VGND VGND VPWR
+ VPWR __dut__._1984_/X sky130_fd_sc_hd__a21o_4
XFILLER_133_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2605_ rst VGND VGND VPWR VPWR __dut__._2605_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2536_ rst VGND VGND VPWR VPWR __dut__._2536_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2467_ rst VGND VGND VPWR VPWR __dut__._2467_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1418_ __dut__._2044_/A1 __dut__._1416_/X __dut__._1417_/X VGND VGND VPWR
+ VPWR __dut__._2660_/D sky130_fd_sc_hd__a21o_4
X__dut__._2398_ rst VGND VGND VPWR VPWR __dut__._2398_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1349_ __dut__._1433_/A __dut__._2642_/Q VGND VGND VPWR VPWR __dut__._1349_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_228_ _297_/Q _227_/B _217_/X VGND VGND VPWR VPWR _300_/D sky130_fd_sc_hd__o21a_4
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_159_ _192_/B VGND VGND VPWR VPWR _171_/B sky130_fd_sc_hd__buf_2
XFILLER_155_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_256_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2249__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1456__A2 mp[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2399__CLK __dut__.__uuf__._2402_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1722_ __dut__.__uuf__._1722_/A VGND VGND VPWR VPWR __dut__._1960_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1653_ __dut__.__uuf__._1654_/A VGND VGND VPWR VPWR __dut__.__uuf__._1653_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2624__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1584_ __dut__.__uuf__._1586_/A VGND VGND VPWR VPWR __dut__.__uuf__._1584_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1392__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2205_ VGND VGND VPWR VPWR __dut__.__uuf__._2205_/HI tie[150] sky130_fd_sc_hd__conb_1
XFILLER_130_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2136_ VGND VGND VPWR VPWR __dut__.__uuf__._2136_/HI tie[81] sky130_fd_sc_hd__conb_1
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2067_ VGND VGND VPWR VPWR __dut__.__uuf__._2067_/HI tie[12] sky130_fd_sc_hd__conb_1
X__dut__._2321_ __dut__._2321_/A __dut__._2321_/B VGND VGND VPWR VPWR __dut__._2321_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2252_ __dut__._2256_/A1 __dut__._2252_/A2 __dut__._2251_/X VGND VGND VPWR
+ VPWR __dut__._2252_/X sky130_fd_sc_hd__a21o_4
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2183_ __dut__._2189_/A __dut__._2183_/B VGND VGND VPWR VPWR __dut__._2183_/X
+ sky130_fd_sc_hd__and2_4
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_127 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1572_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_116 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1534_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_105 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2098_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_138 __dut__._1772_/A1 VGND VGND VPWR VPWR psn_inst_psn_buff_193/A
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_149 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1664_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_149_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2534__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1967_ __dut__._2213_/A __dut__._1967_/B VGND VGND VPWR VPWR __dut__._1967_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1898_ __dut__._1898_/A1 prod[6] __dut__._1897_/X VGND VGND VPWR VPWR __dut__._2868_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2519_ rst VGND VGND VPWR VPWR __dut__._2519_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2444__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2619__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1523__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1155__A __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1705_ __dut__._2347_/B __dut__.__uuf__._1702_/X __dut__._2283_/B
+ __dut__.__uuf__._1703_/X VGND VGND VPWR VPWR prod[26] sky130_fd_sc_hd__o22a_4
XFILLER_119_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2870_ __dut__._2885_/CLK __dut__._2870_/D __dut__._2382_/Y VGND VGND VPWR
+ VPWR __dut__._2870_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1636_ __dut__.__uuf__._1636_/A VGND VGND VPWR VPWR __dut__.__uuf__._1636_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1821_ __dut__._1853_/A __dut__._2829_/Q VGND VGND VPWR VPWR __dut__._1821_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_119_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1567_ __dut__.__uuf__._1564_/X __dut__.__uuf__._1559_/X __dut__._2095_/B
+ __dut__.__uuf__._1548_/X __dut__.__uuf__._1566_/X VGND VGND VPWR VPWR __dut__._2094_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_123_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_5_12_0_tck clkbuf_4_6_0_tck/X VGND VGND VPWR VPWR __dut__._2661_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_134_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1752_ __dut__._1854_/A1 tie[103] __dut__._1751_/X VGND VGND VPWR VPWR __dut__._2795_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1498_ __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR __dut__.__uuf__._1581_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_150_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1683_ __dut__._1701_/A __dut__._2760_/Q VGND VGND VPWR VPWR __dut__._1683_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_130_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_27_0_tck clkbuf_5_27_0_tck/A VGND VGND VPWR VPWR _193_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_48_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2119_ VGND VGND VPWR VPWR __dut__.__uuf__._2119_/HI tie[64] sky130_fd_sc_hd__conb_1
XFILLER_57_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2304_ __dut__._2356_/A1 __dut__._2304_/A2 __dut__._2303_/X VGND VGND VPWR
+ VPWR __dut__._2304_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2529__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2235_ __dut__._2239_/A __dut__._2235_/B VGND VGND VPWR VPWR __dut__._2235_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_60_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2166_ __dut__._2166_/A1 __dut__._2166_/A2 __dut__._2165_/X VGND VGND VPWR
+ VPWR __dut__._2166_/X sky130_fd_sc_hd__a21o_4
X__dut__._2097_ __dut__._2097_/A __dut__._2097_/B VGND VGND VPWR VPWR __dut__._2097_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1356__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2801__CLK clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2439__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1343__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_121_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_219_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1703__A __dut__._1528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1421_ __dut__.__uuf__._1418_/X __dut__.__uuf__._1420_/X __dut__._2161_/B
+ __dut__.__uuf__._1418_/X VGND VGND VPWR VPWR __dut__._2160_/A2 sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._1898__A2 prod[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1352_ __dut__.__uuf__._1351_/Y __dut__.__uuf__._1336_/X __dut__.__uuf__._1337_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1352_/X sky130_fd_sc_hd__o21a_4
XFILLER_131_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1283_ __dut__.__uuf__._1414_/A VGND VGND VPWR VPWR __dut__.__uuf__._1283_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_112_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2020_ __dut__._2024_/A1 __dut__._2020_/A2 __dut__._2019_/X VGND VGND VPWR
+ VPWR __dut__._2020_/X sky130_fd_sc_hd__a21o_4
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1619_ __dut__.__uuf__._1643_/A VGND VGND VPWR VPWR __dut__.__uuf__._1624_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2853_ clkbuf_5_5_0_tck/X __dut__._2853_/D __dut__._2399_/Y VGND VGND VPWR
+ VPWR __dut__._2853_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1804_ __dut__._1804_/A1 tie[129] __dut__._1803_/X VGND VGND VPWR VPWR __dut__._2821_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2784_ __dut__._2885_/CLK __dut__._2784_/D __dut__._2468_/Y VGND VGND VPWR
+ VPWR __dut__._2784_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1735_ __dut__._2327_/A __dut__._2786_/Q VGND VGND VPWR VPWR __dut__._1735_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_89_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1666_ __dut__._1666_/A1 tie[60] __dut__._1665_/X VGND VGND VPWR VPWR __dut__._2752_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1597_ __dut__._1793_/A __dut__._2717_/Q VGND VGND VPWR VPWR __dut__._1597_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2218_ __dut__._2228_/A1 __dut__._2218_/A2 __dut__._2217_/X VGND VGND VPWR
+ VPWR __dut__._2218_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2149_ __dut__._2149_/A __dut__._2149_/B VGND VGND VPWR VPWR __dut__._2149_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_9_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_169_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_336_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1970_ __dut__._2055_/B __dut__._2061_/B __dut__.__uuf__._1969_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1971_/C sky130_fd_sc_hd__o21ai_4
XFILLER_36_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2847__CLK clkbuf_5_4_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1801__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1404_ __dut__.__uuf__._1429_/A VGND VGND VPWR VPWR __dut__.__uuf__._1404_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2384_ __dut__.__uuf__._2422_/CLK __dut__._2272_/X __dut__.__uuf__._1168_/X
+ VGND VGND VPWR VPWR __dut__._2273_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_132_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1335_ __dut__.__uuf__._1771_/A VGND VGND VPWR VPWR __dut__.__uuf__._1711_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_120_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1520_ __dut__._1282_/Y mp[31] __dut__._1519_/X VGND VGND VPWR VPWR __dut__._1520_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_116_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1266_ __dut__._2219_/B __dut__._2217_/B VGND VGND VPWR VPWR __dut__.__uuf__._1266_/X
+ sky130_fd_sc_hd__or2_4
X__dut__.__uuf__._1197_ __dut__.__uuf__._1206_/A VGND VGND VPWR VPWR __dut__.__uuf__._1197_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1451_ _234_/Y __dut__._2669_/Q VGND VGND VPWR VPWR __dut__._1451_/X sky130_fd_sc_hd__and2_4
XFILLER_74_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1382_ __dut__._1382_/A1 __dut__._1380_/X __dut__._1381_/X VGND VGND VPWR
+ VPWR __dut__._2651_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2079__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2003_ __dut__._2213_/A __dut__._2003_/B VGND VGND VPWR VPWR __dut__._2003_/X
+ sky130_fd_sc_hd__and2_4
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_261_ _193_/A _261_/D VGND VGND VPWR VPWR _261_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_psn_inst_psn_buff_22_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_192_ _258_/Q _192_/B VGND VGND VPWR VPWR _257_/D sky130_fd_sc_hd__or2_4
XFILLER_50_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2542__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2836_ __dut__._2845_/CLK __dut__._2836_/D __dut__._2416_/Y VGND VGND VPWR
+ VPWR __dut__._2836_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2767_ __dut__._2767_/CLK __dut__._2767_/D __dut__._2485_/Y VGND VGND VPWR
+ VPWR __dut__._2767_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1718_ __dut__._1726_/A1 tie[86] __dut__._1717_/X VGND VGND VPWR VPWR __dut__._2778_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2698_ __dut__._2721_/CLK __dut__._2698_/D __dut__._2554_/Y VGND VGND VPWR
+ VPWR __dut__._2698_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1649_ __dut__._1661_/A __dut__._2743_/Q VGND VGND VPWR VPWR __dut__._1649_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2282__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_92_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_2_0_tck clkbuf_4_3_0_tck/A VGND VGND VPWR VPWR clkbuf_5_5_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_118_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2452__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_286_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1120_ __dut__.__uuf__._1149_/A VGND VGND VPWR VPWR __dut__.__uuf__._1132_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_102_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1051_ __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR __dut__.__uuf__._1051_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1953_ __dut__.__uuf__._1985_/A __dut__.__uuf__._1953_/B __dut__.__uuf__._1953_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1954_/A sky130_fd_sc_hd__or3_4
XFILLER_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1531__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1884_ __dut__._2023_/B __dut__._2029_/B __dut__.__uuf__._1883_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1885_/C sky130_fd_sc_hd__o21ai_4
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2362__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2621_ rst VGND VGND VPWR VPWR __dut__._2621_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2367_ __dut__.__uuf__._2372_/CLK __dut__._2238_/X __dut__.__uuf__._1217_/X
+ VGND VGND VPWR VPWR __dut__._2239_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2552_ rst VGND VGND VPWR VPWR __dut__._2552_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2298_ __dut__.__uuf__._2319_/CLK __dut__._2100_/X __dut__.__uuf__._1552_/X
+ VGND VGND VPWR VPWR __dut__._2101_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1318_ __dut__.__uuf__._1315_/X __dut__.__uuf__._1317_/X __dut__._2201_/B
+ __dut__.__uuf__._1315_/X VGND VGND VPWR VPWR __dut__._2200_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2483_ rst VGND VGND VPWR VPWR __dut__._2483_/Y sky130_fd_sc_hd__inv_2
X__dut__._1503_ _234_/Y __dut__._2682_/Q VGND VGND VPWR VPWR __dut__._1503_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1249_ __dut__.__uuf__._1249_/A VGND VGND VPWR VPWR __dut__.__uuf__._1249_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1434_ __dut__._1434_/A1 __dut__._1432_/X __dut__._1433_/X VGND VGND VPWR
+ VPWR __dut__._2664_/D sky130_fd_sc_hd__a21o_4
XFILLER_36_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1365_ __dut__._1365_/A __dut__._2646_/Q VGND VGND VPWR VPWR __dut__._1365_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1296_ __dut__._1282_/Y mc[12] __dut__._1295_/X VGND VGND VPWR VPWR __dut__._1296_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2537__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_313_ _193_/A _313_/D trst VGND VGND VPWR VPWR _313_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_244_ _202_/X _293_/Q VGND VGND VPWR VPWR _244_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_175_ _182_/A VGND VGND VPWR VPWR _181_/B sky130_fd_sc_hd__buf_2
XFILLER_155_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1704__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2819_ clkbuf_5_1_0_tck/X __dut__._2819_/D __dut__._2433_/Y VGND VGND VPWR
+ VPWR __dut__._2819_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_111_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2692__CLK clkbuf_5_2_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2447__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1351__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1711__A __dut__.__uuf__._1711_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2221_ VGND VGND VPWR VPWR __dut__.__uuf__._2221_/HI tie[166] sky130_fd_sc_hd__conb_1
XFILLER_88_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2152_ VGND VGND VPWR VPWR __dut__.__uuf__._2152_/HI tie[97] sky130_fd_sc_hd__conb_1
XFILLER_102_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2083_ VGND VGND VPWR VPWR __dut__.__uuf__._2083_/HI tie[28] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1103_ __dut__.__uuf__._1103_/A VGND VGND VPWR VPWR __dut__.__uuf__._1103_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_84_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1034_ __dut__.__uuf__._1103_/A VGND VGND VPWR VPWR __dut__.__uuf__._1034_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_84_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2357__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_309 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1293_/A
+ sky130_fd_sc_hd__buf_2
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1936_ __dut__._2043_/B __dut__._2049_/B VGND VGND VPWR VPWR __dut__.__uuf__._1937_/A
+ sky130_fd_sc_hd__and2_4
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1867_ __dut__.__uuf__._1867_/A VGND VGND VPWR VPWR __dut__._2016_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1046__B2 __dut__.__uuf__._1040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1798_ __dut__.__uuf__._1798_/A __dut__.__uuf__._1798_/B __dut__.__uuf__._1798_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1799_/A sky130_fd_sc_hd__or3_4
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1983_ __dut__._2213_/A __dut__._1983_/B VGND VGND VPWR VPWR __dut__._1983_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2419_ __dut__.__uuf__._2422_/CLK __dut__._2342_/X __dut__.__uuf__._1063_/X
+ VGND VGND VPWR VPWR __dut__._2343_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_154_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2604_ rst VGND VGND VPWR VPWR __dut__._2604_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0___dut__.__uuf__.__clk_source__ clkbuf_2_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
X__dut__._2535_ rst VGND VGND VPWR VPWR __dut__._2535_/Y sky130_fd_sc_hd__inv_2
X__dut__._2466_ rst VGND VGND VPWR VPWR __dut__._2466_/Y sky130_fd_sc_hd__inv_2
X__dut__._2397_ rst VGND VGND VPWR VPWR __dut__._2397_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1417_ __dut__._1417_/A __dut__._2649_/Q VGND VGND VPWR VPWR __dut__._1417_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1348_ __dut__._1282_/Y mc[24] __dut__._1347_/X VGND VGND VPWR VPWR __dut__._1348_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2320__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0___dut__.__uuf__.__clk_source___A clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_227_ _231_/A _227_/B VGND VGND VPWR VPWR _299_/D sky130_fd_sc_hd__and2_4
XFILLER_156_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_158_ _287_/Q _163_/B VGND VGND VPWR VPWR _286_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2350__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__239__A1 tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_249_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_151_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1721_ __dut__.__uuf__._1768_/A __dut__.__uuf__._1721_/B __dut__.__uuf__._1721_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1722_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1652_ __dut__.__uuf__._1654_/A VGND VGND VPWR VPWR __dut__.__uuf__._1652_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_21_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1583_ __dut__.__uuf__._1586_/A VGND VGND VPWR VPWR __dut__.__uuf__._1583_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_134_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1392__A2 mp[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2204_ VGND VGND VPWR VPWR __dut__.__uuf__._2204_/HI tie[149] sky130_fd_sc_hd__conb_1
XFILLER_115_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2135_ VGND VGND VPWR VPWR __dut__.__uuf__._2135_/HI tie[80] sky130_fd_sc_hd__conb_1
XFILLER_124_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2066_ VGND VGND VPWR VPWR __dut__.__uuf__._2066_/HI tie[11] sky130_fd_sc_hd__conb_1
X__dut__._2320_ __dut__._2322_/A1 __dut__._2320_/A2 __dut__._2319_/X VGND VGND VPWR
+ VPWR __dut__._2320_/X sky130_fd_sc_hd__a21o_4
X__dut__._2251_ __dut__._2251_/A __dut__._2251_/B VGND VGND VPWR VPWR __dut__._2251_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2087__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2182_ __dut__._2182_/A1 __dut__._2182_/A2 __dut__._2181_/X VGND VGND VPWR
+ VPWR __dut__._2182_/X sky130_fd_sc_hd__a21o_4
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_128 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1570_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_117 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1538_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_106 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._2096_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_33_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_139 psn_inst_psn_buff_193/A VGND VGND VPWR VPWR __dut__._1494_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1919_ __dut__.__uuf__._1875_/X __dut__.__uuf__._1917_/B __dut__.__uuf__._1917_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1920_/C sky130_fd_sc_hd__o21a_4
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1966_ __dut__._2078_/A1 __dut__._1966_/A2 __dut__._1965_/X VGND VGND VPWR
+ VPWR __dut__._1966_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2550__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1897_ __dut__._1897_/A __dut__._2867_/Q VGND VGND VPWR VPWR __dut__._1897_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_4_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2518_ rst VGND VGND VPWR VPWR __dut__._2518_/Y sky130_fd_sc_hd__inv_2
X__dut__._2449_ rst VGND VGND VPWR VPWR __dut__._2449_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2460__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1704_ __dut__._2345_/B __dut__.__uuf__._1702_/X __dut__._2281_/B
+ __dut__.__uuf__._1703_/X VGND VGND VPWR VPWR prod[25] sky130_fd_sc_hd__o22a_4
XANTENNA___dut__.__uuf__._1171__A __dut__.__uuf__._1215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1635_ __dut__.__uuf__._1636_/A VGND VGND VPWR VPWR __dut__.__uuf__._1635_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1820_ __dut__._1854_/A1 tie[137] __dut__._1819_/X VGND VGND VPWR VPWR __dut__._2829_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_119_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1566_ __dut__._1400_/X __dut__.__uuf__._1565_/X __dut__._2097_/B
+ __dut__.__uuf__._1549_/X VGND VGND VPWR VPWR __dut__.__uuf__._1566_/X sky130_fd_sc_hd__o22a_4
XFILLER_150_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1751_ __dut__._1853_/A __dut__._2794_/Q VGND VGND VPWR VPWR __dut__._1751_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2370__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1497_ __dut__.__uuf__._1478_/X __dut__.__uuf__._1495_/X __dut__._2127_/B
+ __dut__.__uuf__._1484_/X __dut__.__uuf__._1496_/X VGND VGND VPWR VPWR __dut__._2126_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_135_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1682_ __dut__._1682_/A1 tie[68] __dut__._1681_/X VGND VGND VPWR VPWR __dut__._2760_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2118_ VGND VGND VPWR VPWR __dut__.__uuf__._2118_/HI tie[63] sky130_fd_sc_hd__conb_1
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2303_ __dut__._2313_/A __dut__._2303_/B VGND VGND VPWR VPWR __dut__._2303_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._2049_ __dut__.__uuf__._2042_/A __dut__.__uuf__._2047_/B __dut__.__uuf__._1038_/X
+ VGND VGND VPWR VPWR __dut__._2082_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2234_ __dut__._2356_/A1 __dut__._2234_/A2 __dut__._2233_/X VGND VGND VPWR
+ VPWR __dut__._2234_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_52_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2165_ __dut__._2167_/A __dut__._2165_/B VGND VGND VPWR VPWR __dut__._2165_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2545__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2096_ __dut__._2096_/A1 __dut__._2096_/A2 __dut__._2095_/X VGND VGND VPWR
+ VPWR __dut__._2096_/X sky130_fd_sc_hd__a21o_4
XFILLER_60_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2239__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_138_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1356__A2 mc[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1949_ __dut__._1949_/A __dut__._2893_/Q VGND VGND VPWR VPWR __dut__._1949_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1292__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_psn_inst_psn_buff_114_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2455__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1420_ __dut__.__uuf__._1419_/Y __dut__.__uuf__._1413_/X __dut__.__uuf__._1414_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1420_/X sky130_fd_sc_hd__o21a_4
XFILLER_156_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1351_ __dut__._2189_/B VGND VGND VPWR VPWR __dut__.__uuf__._1351_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_132_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1282_ __dut__._1520_/X __dut__.__uuf__._1307_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1414_/A sky130_fd_sc_hd__nand2_4
XFILLER_131_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2365__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1618_ __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR __dut__.__uuf__._1643_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._2852_ clkbuf_5_6_0_tck/X __dut__._2852_/D __dut__._2400_/Y VGND VGND VPWR
+ VPWR __dut__._2852_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1803_ __dut__._2213_/A __dut__._2820_/Q VGND VGND VPWR VPWR __dut__._1803_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2783_ __dut__._2885_/CLK __dut__._2783_/D __dut__._2469_/Y VGND VGND VPWR
+ VPWR __dut__._2783_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1549_ __dut__.__uuf__._1771_/A VGND VGND VPWR VPWR __dut__.__uuf__._1549_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1734_ __dut__._1910_/A1 tie[94] __dut__._1733_/X VGND VGND VPWR VPWR __dut__._2786_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_89_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1665_ __dut__._1665_/A __dut__._2751_/Q VGND VGND VPWR VPWR __dut__._1665_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1596_ __dut__._1790_/A1 tie[25] __dut__._1595_/X VGND VGND VPWR VPWR __dut__._2717_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2217_ __dut__._2217_/A __dut__._2217_/B VGND VGND VPWR VPWR __dut__._2217_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2649__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2148_ __dut__._2228_/A1 __dut__._2148_/A2 __dut__._2147_/X VGND VGND VPWR
+ VPWR __dut__._2148_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2079_ __dut__._2213_/A __dut__._2079_/B VGND VGND VPWR VPWR __dut__._2079_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_126_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2799__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_329_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_231_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_11_0_tck clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR __dut__._2357_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_26_0_tck clkbuf_5_27_0_tck/A VGND VGND VPWR VPWR _312_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2383_ __dut__.__uuf__._2415_/CLK __dut__._2270_/X __dut__.__uuf__._1170_/X
+ VGND VGND VPWR VPWR __dut__._2271_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1403_ __dut__.__uuf__._1402_/Y __dut__.__uuf__._1388_/X __dut__.__uuf__._1389_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1403_/X sky130_fd_sc_hd__o21a_4
XFILLER_132_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1334_ __dut__._2195_/B VGND VGND VPWR VPWR __dut__.__uuf__._1334_/Y
+ sky130_fd_sc_hd__inv_2
Xclkbuf_4_3_0___dut__.__uuf__.__clk_source__ clkbuf_4_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2323_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1265_ __dut__.__uuf__._1269_/A VGND VGND VPWR VPWR __dut__.__uuf__._1265_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_58_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1450_ __dut__._1450_/A1 __dut__._1448_/X __dut__._1449_/X VGND VGND VPWR
+ VPWR __dut__._2668_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1196_ __dut__.__uuf__._1192_/X __dut__.__uuf__._1188_/X __dut__._2255_/B
+ __dut__._2257_/B __dut__.__uuf__._1185_/X VGND VGND VPWR VPWR __dut__._2254_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_132_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1381_ __dut__._2095_/A __dut__._2650_/Q VGND VGND VPWR VPWR __dut__._1381_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_27_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2002_ __dut__._2008_/A1 __dut__._2002_/A2 __dut__._2001_/X VGND VGND VPWR
+ VPWR __dut__._2002_/X sky130_fd_sc_hd__a21o_4
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_260_ _193_/A _260_/D VGND VGND VPWR VPWR _260_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_191_ _259_/Q _192_/B VGND VGND VPWR VPWR _258_/D sky130_fd_sc_hd__or2_4
XFILLER_41_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_psn_inst_psn_buff_15_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2835_ __dut__._2845_/CLK __dut__._2835_/D __dut__._2417_/Y VGND VGND VPWR
+ VPWR __dut__._2835_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1439__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2766_ __dut__._2865_/CLK __dut__._2766_/D __dut__._2486_/Y VGND VGND VPWR
+ VPWR __dut__._2766_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1717_ __dut__._1729_/A __dut__._2777_/Q VGND VGND VPWR VPWR __dut__._1717_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2697_ __dut__._2721_/CLK __dut__._2697_/D __dut__._2555_/Y VGND VGND VPWR
+ VPWR __dut__._2697_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1648_ __dut__._1658_/A1 tie[51] __dut__._1647_/X VGND VGND VPWR VPWR __dut__._2743_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1579_ __dut__._1793_/A __dut__._2708_/Q VGND VGND VPWR VPWR __dut__._1579_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_181_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_279_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1050_ __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR __dut__.__uuf__._1229_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1952_ __dut__.__uuf__._1929_/X __dut__.__uuf__._1950_/B __dut__.__uuf__._1950_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1953_/C sky130_fd_sc_hd__o21a_4
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1883_ __dut__.__uuf__._1883_/A VGND VGND VPWR VPWR __dut__.__uuf__._1883_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2620_ rst VGND VGND VPWR VPWR __dut__._2620_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2366_ __dut__.__uuf__._2372_/CLK __dut__._2236_/X __dut__.__uuf__._1220_/X
+ VGND VGND VPWR VPWR __dut__._2237_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_132_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2551_ rst VGND VGND VPWR VPWR __dut__._2551_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2297_ __dut__.__uuf__._2319_/CLK __dut__._2098_/X __dut__.__uuf__._1555_/X
+ VGND VGND VPWR VPWR __dut__._2099_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1317_ __dut__.__uuf__._1316_/Y __dut__.__uuf__._1309_/X __dut__.__uuf__._1311_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1317_/X sky130_fd_sc_hd__o21a_4
XFILLER_98_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1502_ __dut__._1616_/A1 __dut__._1500_/X __dut__._1501_/X VGND VGND VPWR
+ VPWR __dut__._2681_/D sky130_fd_sc_hd__a21o_4
X__dut__._2482_ rst VGND VGND VPWR VPWR __dut__._2482_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1248_ __dut__.__uuf__._1229_/A __dut__.__uuf__._1241_/X __dut__.__uuf__._1242_/X
+ __dut__._2229_/B __dut__.__uuf__._1247_/X VGND VGND VPWR VPWR __dut__._2228_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_47_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1433_ __dut__._1433_/A __dut__._2663_/Q VGND VGND VPWR VPWR __dut__._1433_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1179_ __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR __dut__.__uuf__._1190_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_101_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1364_ __dut__._1282_/Y mc[28] __dut__._1363_/X VGND VGND VPWR VPWR __dut__._1364_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1295_ _234_/Y __dut__._2630_/Q VGND VGND VPWR VPWR __dut__._1295_/X sky130_fd_sc_hd__and2_4
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ _312_/CLK _312_/D trst VGND VGND VPWR VPWR _312_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_243_ tdi _153_/C _300_/Q _313_/Q VGND VGND VPWR VPWR _313_/D sky130_fd_sc_hd__o22a_4
XFILLER_156_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2553__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_174_ _274_/Q _186_/B VGND VGND VPWR VPWR _273_/D sky130_fd_sc_hd__or2_4
XFILLER_155_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0___dut__.__uuf__.__clk_source___A clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2818_ clkbuf_5_0_0_tck/X __dut__._2818_/D __dut__._2434_/Y VGND VGND VPWR
+ VPWR __dut__._2818_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2837__CLK __dut__._2845_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2749_ __dut__._2894_/CLK __dut__._2749_/D __dut__._2503_/Y VGND VGND VPWR
+ VPWR __dut__._2749_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1468__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2463__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2220_ VGND VGND VPWR VPWR __dut__.__uuf__._2220_/HI tie[165] sky130_fd_sc_hd__conb_1
XFILLER_115_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1807__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2151_ VGND VGND VPWR VPWR __dut__.__uuf__._2151_/HI tie[96] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2082_ VGND VGND VPWR VPWR __dut__.__uuf__._2082_/HI tie[27] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1102_ __dut__.__uuf__._1102_/A VGND VGND VPWR VPWR __dut__.__uuf__._1102_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_84_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1033_ __dut__.__uuf__._1564_/A VGND VGND VPWR VPWR __dut__.__uuf__._1103_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_110_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1935_ __dut__._1332_/X VGND VGND VPWR VPWR __dut__.__uuf__._1939_/B
+ sky130_fd_sc_hd__inv_2
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1866_ __dut__.__uuf__._1877_/A __dut__.__uuf__._1866_/B __dut__.__uuf__._1866_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1867_/A sky130_fd_sc_hd__or3_4
XANTENNA___dut__.__uuf__._1046__A2 __dut__.__uuf__._1038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2373__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1797_ __dut__._1991_/B __dut__._1997_/B __dut__.__uuf__._1796_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1798_/C sky130_fd_sc_hd__o21ai_4
XFILLER_149_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1934__A2 prod[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1982_ __dut__._2000_/A1 __dut__._1982_/A2 __dut__._1981_/X VGND VGND VPWR
+ VPWR __dut__._1982_/X sky130_fd_sc_hd__a21o_4
XFILLER_152_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1698__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2418_ __dut__.__uuf__._2422_/CLK __dut__._2340_/X __dut__.__uuf__._1065_/X
+ VGND VGND VPWR VPWR __dut__._2341_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2603_ rst VGND VGND VPWR VPWR __dut__._2603_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2349_ __dut__.__uuf__._2355_/CLK __dut__._2202_/X __dut__.__uuf__._1305_/X
+ VGND VGND VPWR VPWR __dut__._2203_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_121_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2534_ rst VGND VGND VPWR VPWR __dut__._2534_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_1_0_tck clkbuf_4_1_0_tck/A VGND VGND VPWR VPWR clkbuf_5_3_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_87_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_82_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2465_ rst VGND VGND VPWR VPWR __dut__._2465_/Y sky130_fd_sc_hd__inv_2
X__dut__._2396_ rst VGND VGND VPWR VPWR __dut__._2396_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2548__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1416_ __dut__._1282_/Y mc[3] __dut__._1415_/X VGND VGND VPWR VPWR __dut__._1416_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1347_ _234_/Y __dut__._2643_/Q VGND VGND VPWR VPWR __dut__._1347_/X sky130_fd_sc_hd__and2_4
XFILLER_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_226_ _300_/Q _301_/Q VGND VGND VPWR VPWR _227_/B sky130_fd_sc_hd__or2_4
X_157_ _288_/Q _163_/B VGND VGND VPWR VPWR _287_/D sky130_fd_sc_hd__and2_4
XFILLER_112_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2458__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_144_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_311_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1720_ __dut__.__uuf__._1276_/X __dut__.__uuf__._1718_/B __dut__.__uuf__._1718_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1721_/C sky130_fd_sc_hd__o21a_4
XFILLER_147_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1651_ __dut__.__uuf__._1654_/A VGND VGND VPWR VPWR __dut__.__uuf__._1651_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2295__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2193__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1582_ __dut__.__uuf__._1586_/A VGND VGND VPWR VPWR __dut__.__uuf__._1582_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_134_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2203_ VGND VGND VPWR VPWR __dut__.__uuf__._2203_/HI tie[148] sky130_fd_sc_hd__conb_1
XFILLER_115_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2134_ VGND VGND VPWR VPWR __dut__.__uuf__._2134_/HI tie[79] sky130_fd_sc_hd__conb_1
XFILLER_69_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2065_ VGND VGND VPWR VPWR __dut__.__uuf__._2065_/HI tie[10] sky130_fd_sc_hd__conb_1
XFILLER_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2368__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2250_ __dut__._2256_/A1 __dut__._2250_/A2 __dut__._2249_/X VGND VGND VPWR
+ VPWR __dut__._2250_/X sky130_fd_sc_hd__a21o_4
XFILLER_29_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1852__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2181_ __dut__._2189_/A __dut__._2181_/B VGND VGND VPWR VPWR __dut__._2181_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_140_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_118 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1542_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_107 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1366_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_129 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1568_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1918_ __dut__.__uuf__._1918_/A VGND VGND VPWR VPWR __dut__.__uuf__._1920_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_24_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1849_ __dut__._2011_/B __dut__._2017_/B VGND VGND VPWR VPWR __dut__.__uuf__._1850_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2682__CLK clkbuf_5_3_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1965_ __dut__._2213_/A __dut__._1965_/B VGND VGND VPWR VPWR __dut__._1965_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_79_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1447__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1896_ __dut__._1896_/A1 prod[5] __dut__._1895_/X VGND VGND VPWR VPWR __dut__._2867_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_59_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2517_ rst VGND VGND VPWR VPWR __dut__._2517_/Y sky130_fd_sc_hd__inv_2
X__dut__._2448_ rst VGND VGND VPWR VPWR __dut__._2448_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2379_ rst VGND VGND VPWR VPWR __dut__._2379_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_209_ _208_/Y _209_/A2 _245_/Q _251_/Q VGND VGND VPWR VPWR _210_/B sky130_fd_sc_hd__o22a_4
XFILLER_143_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_261_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1834__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1703_ __dut__._1528_/X VGND VGND VPWR VPWR __dut__.__uuf__._1703_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1634_ __dut__.__uuf__._1636_/A VGND VGND VPWR VPWR __dut__.__uuf__._1634_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_119_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1565_ __dut__.__uuf__._1565_/A VGND VGND VPWR VPWR __dut__.__uuf__._1565_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1750_ __dut__._1854_/A1 tie[102] __dut__._1749_/X VGND VGND VPWR VPWR __dut__._2794_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2801__D __dut__._2801_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._1496_ __dut__._1472_/X __dut__.__uuf__._1480_/X __dut__._2129_/B
+ __dut__.__uuf__._1485_/X VGND VGND VPWR VPWR __dut__.__uuf__._1496_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1681_ __dut__._1701_/A __dut__._2759_/Q VGND VGND VPWR VPWR __dut__._1681_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2310__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_142_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2117_ VGND VGND VPWR VPWR __dut__.__uuf__._2117_/HI tie[62] sky130_fd_sc_hd__conb_1
X__dut__._2302_ __dut__._2356_/A1 __dut__._2302_/A2 __dut__._2301_/X VGND VGND VPWR
+ VPWR __dut__._2302_/X sky130_fd_sc_hd__a21o_4
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2048_ __dut__.__uuf__._2048_/A VGND VGND VPWR VPWR __dut__._2084_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_84_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2233_ __dut__._2313_/A __dut__._2233_/B VGND VGND VPWR VPWR __dut__._2233_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_72_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2164_ __dut__._2166_/A1 __dut__._2164_/A2 __dut__._2163_/X VGND VGND VPWR
+ VPWR __dut__._2164_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_45_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2095_ __dut__._2095_/A __dut__._2095_/B VGND VGND VPWR VPWR __dut__._2095_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1362__A __dut__.__uuf__._1711_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2561__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1948_ __dut__._2328_/A1 prod[31] __dut__._1947_/X VGND VGND VPWR VPWR __dut__._2893_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1879_ __dut__._2213_/A __dut__._2858_/Q VGND VGND VPWR VPWR __dut__._1879_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__271__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1816__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1292__A2 mc[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__156__A tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_107_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2471__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1350_ __dut__.__uuf__._1350_/A VGND VGND VPWR VPWR __dut__.__uuf__._1350_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_132_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1281_ __dut__._2213_/B VGND VGND VPWR VPWR __dut__.__uuf__._1281_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_124_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2232__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2851_ clkbuf_5_6_0_tck/X __dut__._2851_/D __dut__._2401_/Y VGND VGND VPWR
+ VPWR __dut__._2851_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2381__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1617_ __dut__.__uuf__._1617_/A VGND VGND VPWR VPWR __dut__.__uuf__._1617_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1802_ __dut__._1802_/A1 tie[128] __dut__._1801_/X VGND VGND VPWR VPWR __dut__._2820_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2782_ __dut__._2885_/CLK __dut__._2782_/D __dut__._2470_/Y VGND VGND VPWR
+ VPWR __dut__._2782_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1548_ __dut__.__uuf__._1548_/A VGND VGND VPWR VPWR __dut__.__uuf__._1548_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1733_ __dut__._1733_/A __dut__._2785_/Q VGND VGND VPWR VPWR __dut__._1733_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1479_ __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR __dut__.__uuf__._1565_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_103_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1664_ __dut__._1664_/A1 tie[59] __dut__._1663_/X VGND VGND VPWR VPWR __dut__._2751_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_131_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1595_ __dut__._1793_/A __dut__._2716_/Q VGND VGND VPWR VPWR __dut__._1595_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2216_ __dut__._2228_/A1 __dut__._2216_/A2 __dut__._2215_/X VGND VGND VPWR
+ VPWR __dut__._2216_/X sky130_fd_sc_hd__a21o_4
XFILLER_33_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2556__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2147_ __dut__._2147_/A __dut__._2147_/B VGND VGND VPWR VPWR __dut__._2147_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2078_ __dut__._2078_/A1 __dut__._2078_/A2 __dut__._2077_/X VGND VGND VPWR
+ VPWR __dut__._2078_/X sky130_fd_sc_hd__a21o_4
XFILLER_145_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2291__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2466__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_290 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2107_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_145_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1402_ __dut__._2169_/B VGND VGND VPWR VPWR __dut__.__uuf__._1402_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_144_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2382_ __dut__.__uuf__._2415_/CLK __dut__._2268_/X __dut__.__uuf__._1173_/X
+ VGND VGND VPWR VPWR __dut__._2269_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_104_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1333_ __dut__.__uuf__._1350_/A VGND VGND VPWR VPWR __dut__.__uuf__._1333_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1264_ __dut__.__uuf__._1236_/A __dut__.__uuf__._1263_/Y __dut__.__uuf__._1229_/X
+ __dut__._2221_/B __dut__.__uuf__._1247_/X VGND VGND VPWR VPWR __dut__._2220_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_113_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1195_ __dut__.__uuf__._1206_/A VGND VGND VPWR VPWR __dut__.__uuf__._1195_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1177__A __dut__.__uuf__._1177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1380_ __dut__._1282_/Y mc[31] __dut__._1379_/X VGND VGND VPWR VPWR __dut__._1380_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2229__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_82_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2376__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1280__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2001_ __dut__._2213_/A __dut__._2001_/B VGND VGND VPWR VPWR __dut__._2001_/X
+ sky130_fd_sc_hd__and2_4
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_190_ _260_/Q _190_/B VGND VGND VPWR VPWR _259_/D sky130_fd_sc_hd__and2_4
XFILLER_127_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2834_ __dut__._2845_/CLK __dut__._2834_/D __dut__._2418_/Y VGND VGND VPWR
+ VPWR __dut__._2834_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2765_ __dut__._2865_/CLK __dut__._2765_/D __dut__._2487_/Y VGND VGND VPWR
+ VPWR __dut__._2765_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1716_ __dut__._1726_/A1 tie[85] __dut__._1715_/X VGND VGND VPWR VPWR __dut__._2777_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_150_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2696_ clkbuf_5_2_0_tck/X __dut__._2696_/D __dut__._2556_/Y VGND VGND VPWR
+ VPWR __dut__._2696_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1455__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1647_ __dut__._1661_/A __dut__._2742_/Q VGND VGND VPWR VPWR __dut__._1647_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_66_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1578_ __dut__._1578_/A1 tie[16] __dut__._1577_/X VGND VGND VPWR VPWR __dut__._2708_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_64_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_13_0___dut__.__uuf__.__clk_source__ clkbuf_3_6_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2335_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_122_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0___dut__.__uuf__.__clk_source__ __dut__._2358_/X VGND VGND VPWR VPWR clkbuf_0___dut__.__uuf__.__clk_source__/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_174_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1951_ __dut__.__uuf__._1951_/A VGND VGND VPWR VPWR __dut__.__uuf__._1953_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1882_ __dut__._2023_/B __dut__._2029_/B VGND VGND VPWR VPWR __dut__.__uuf__._1883_/A
+ sky130_fd_sc_hd__and2_4
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2365_ __dut__.__uuf__._2372_/CLK __dut__._2234_/X __dut__.__uuf__._1224_/X
+ VGND VGND VPWR VPWR __dut__._2235_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1316_ __dut__._2203_/B VGND VGND VPWR VPWR __dut__.__uuf__._1316_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_132_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2550_ rst VGND VGND VPWR VPWR __dut__._2550_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2296_ __dut__.__uuf__._2319_/CLK __dut__._2096_/X __dut__.__uuf__._1558_/X
+ VGND VGND VPWR VPWR __dut__._2097_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_143_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2481_ rst VGND VGND VPWR VPWR __dut__._2481_/Y sky130_fd_sc_hd__inv_2
X__dut__._1501_ __dut__._1617_/A __dut__._2680_/Q VGND VGND VPWR VPWR __dut__._1501_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1247_ __dut__.__uuf__._1429_/A VGND VGND VPWR VPWR __dut__.__uuf__._1247_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1432_ __dut__._1282_/Y mp[11] __dut__._1431_/X VGND VGND VPWR VPWR __dut__._1432_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1178_ __dut__.__uuf__._1177_/X __dut__.__uuf__._1174_/X __dut__._2267_/B
+ __dut__._2269_/B __dut__.__uuf__._1171_/X VGND VGND VPWR VPWR __dut__._2266_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1363_ _234_/Y __dut__._2647_/Q VGND VGND VPWR VPWR __dut__._1363_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2789__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1294_ __dut__._1564_/A1 __dut__._1292_/X __dut__._1293_/X VGND VGND VPWR
+ VPWR __dut__._2629_/D sky130_fd_sc_hd__a21o_4
XFILLER_15_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__238__B _304_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_311_ _312_/CLK _311_/D trst VGND VGND VPWR VPWR _311_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_156_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_242_ _310_/Q _309_/Q _242_/C _242_/D VGND VGND VPWR VPWR _242_/X sky130_fd_sc_hd__and4_4
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_173_ _192_/B VGND VGND VPWR VPWR _186_/B sky130_fd_sc_hd__buf_2
XFILLER_109_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_10_0_tck clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR __dut__._2721_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2817_ clkbuf_5_0_0_tck/X __dut__._2817_/D __dut__._2435_/Y VGND VGND VPWR
+ VPWR __dut__._2817_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2748_ __dut__._2894_/CLK __dut__._2748_/D __dut__._2504_/Y VGND VGND VPWR
+ VPWR __dut__._2748_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2679_ __dut__._2680_/CLK __dut__._2679_/D __dut__._2573_/Y VGND VGND VPWR
+ VPWR __dut__._2679_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_25_0_tck clkbuf_5_25_0_tck/A VGND VGND VPWR VPWR _288_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1468__A2 mp[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1913__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_291_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2150_ VGND VGND VPWR VPWR __dut__.__uuf__._2150_/HI tie[95] sky130_fd_sc_hd__conb_1
XFILLER_114_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2081_ VGND VGND VPWR VPWR __dut__.__uuf__._2081_/HI tie[26] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._1101_ __dut__.__uuf__._1087_/X __dut__.__uuf__._1100_/X __dut__._2319_/B
+ __dut__._2321_/B __dut__.__uuf__._1097_/X VGND VGND VPWR VPWR __dut__._2318_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1032_ __dut__.__uuf__._1191_/A VGND VGND VPWR VPWR __dut__.__uuf__._1564_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1823__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1455__A __dut__.__uuf__._1478_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1934_ __dut__.__uuf__._1988_/A VGND VGND VPWR VPWR __dut__.__uuf__._1985_/A
+ sky130_fd_sc_hd__buf_2
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1865_ __dut__.__uuf__._1821_/X __dut__.__uuf__._1863_/B __dut__.__uuf__._1863_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1866_/C sky130_fd_sc_hd__o21a_4
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1796_ __dut__.__uuf__._1796_/A VGND VGND VPWR VPWR __dut__.__uuf__._1796_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_149_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1981_ __dut__._2213_/A __dut__._1981_/B VGND VGND VPWR VPWR __dut__._1981_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_138_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2417_ __dut__.__uuf__._2422_/CLK __dut__._2338_/X __dut__.__uuf__._1068_/X
+ VGND VGND VPWR VPWR __dut__._2339_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2602_ rst VGND VGND VPWR VPWR __dut__._2602_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2348_ __dut__.__uuf__._2348_/CLK __dut__._2200_/X __dut__.__uuf__._1314_/X
+ VGND VGND VPWR VPWR __dut__._2201_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2533_ rst VGND VGND VPWR VPWR __dut__._2533_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2279_ __dut__.__uuf__._2288_/CLK __dut__._2062_/X __dut__.__uuf__._1596_/X
+ VGND VGND VPWR VPWR __dut__._2063_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_59_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2464_ rst VGND VGND VPWR VPWR __dut__._2464_/Y sky130_fd_sc_hd__inv_2
X__dut__._2395_ rst VGND VGND VPWR VPWR __dut__._2395_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1415_ _234_/Y __dut__._2660_/Q VGND VGND VPWR VPWR __dut__._1415_/X sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_75_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1346_ __dut__._1346_/A1 __dut__._1344_/X __dut__._1345_/X VGND VGND VPWR
+ VPWR __dut__._2642_/D sky130_fd_sc_hd__a21o_4
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2564__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_225_ _299_/Q _298_/Q _217_/X VGND VGND VPWR VPWR _298_/D sky130_fd_sc_hd__o21a_4
XFILLER_7_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2804__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_156_ tdi _163_/B VGND VGND VPWR VPWR _288_/D sky130_fd_sc_hd__and2_4
XFILLER_124_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_137_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2474__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_304_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1650_ __dut__.__uuf__._1654_/A VGND VGND VPWR VPWR __dut__.__uuf__._1650_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1581_ __dut__.__uuf__._1581_/A VGND VGND VPWR VPWR __dut__.__uuf__._1586_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_146_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2202_ VGND VGND VPWR VPWR __dut__.__uuf__._2202_/HI tie[147] sky130_fd_sc_hd__conb_1
XFILLER_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2133_ VGND VGND VPWR VPWR __dut__.__uuf__._2133_/HI tie[78] sky130_fd_sc_hd__conb_1
XFILLER_130_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2064_ VGND VGND VPWR VPWR __dut__.__uuf__._2064_/HI tie[9] sky130_fd_sc_hd__conb_1
XFILLER_29_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1185__A __dut__.__uuf__._1215_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2180_ __dut__._2180_/A1 __dut__._2180_/A2 __dut__._2179_/X VGND VGND VPWR
+ VPWR __dut__._2180_/X sky130_fd_sc_hd__a21o_4
XFILLER_25_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_119 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1564_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_108 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1462_/A1
+ sky130_fd_sc_hd__buf_2
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__297__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2384__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1917_ __dut__.__uuf__._1960_/A __dut__.__uuf__._1917_/B __dut__.__uuf__._1917_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1918_/A sky130_fd_sc_hd__or3_4
XFILLER_33_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1848_ __dut__._1296_/X VGND VGND VPWR VPWR __dut__.__uuf__._1852_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2827__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1368__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1779_ __dut__.__uuf__._1766_/X __dut__.__uuf__._1777_/B __dut__.__uuf__._1777_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1780_/C sky130_fd_sc_hd__o21a_4
XFILLER_125_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1964_ __dut__._1964_/A1 __dut__._1964_/A2 __dut__._1963_/X VGND VGND VPWR
+ VPWR __dut__._1964_/X sky130_fd_sc_hd__a21o_4
XFILLER_153_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1895_ __dut__._2243_/A __dut__._2866_/Q VGND VGND VPWR VPWR __dut__._1895_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1540__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2516_ rst VGND VGND VPWR VPWR __dut__._2516_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._2559__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2447_ rst VGND VGND VPWR VPWR __dut__._2447_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_9_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1463__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2378_ rst VGND VGND VPWR VPWR __dut__._2378_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1329_ __dut__._2095_/A __dut__._2627_/Q VGND VGND VPWR VPWR __dut__._1329_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_208_ _245_/Q VGND VGND VPWR VPWR _208_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_139_ _139_/A VGND VGND VPWR VPWR _309_/D sky130_fd_sc_hd__inv_2
XFILLER_124_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_254_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2469__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1702_ __dut__.__uuf__._1702_/A VGND VGND VPWR VPWR __dut__.__uuf__._1702_/X
+ sky130_fd_sc_hd__buf_2
Xclkbuf_4_0_0_tck clkbuf_4_1_0_tck/A VGND VGND VPWR VPWR clkbuf_5_1_0_tck/A sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1633_ __dut__.__uuf__._1636_/A VGND VGND VPWR VPWR __dut__.__uuf__._1633_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1564_ __dut__.__uuf__._1564_/A VGND VGND VPWR VPWR __dut__.__uuf__._1564_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1495_ __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR __dut__.__uuf__._1495_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1680_ __dut__._1726_/A1 tie[67] __dut__._1679_/X VGND VGND VPWR VPWR __dut__._2759_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2116_ VGND VGND VPWR VPWR __dut__.__uuf__._2116_/HI tie[61] sky130_fd_sc_hd__conb_1
XANTENNA___dut__._2379__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2301_ __dut__._2313_/A __dut__._2301_/B VGND VGND VPWR VPWR __dut__._2301_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2047_ __dut__.__uuf__._2047_/A __dut__.__uuf__._2047_/B __dut__.__uuf__._2047_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2048_/A sky130_fd_sc_hd__or3_4
X__dut__._2232_ __dut__._2356_/A1 __dut__._2232_/A2 __dut__._2231_/X VGND VGND VPWR
+ VPWR __dut__._2232_/X sky130_fd_sc_hd__a21o_4
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1286__B1 __dut__._1285_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2163_ __dut__._2167_/A __dut__._2163_/B VGND VGND VPWR VPWR __dut__._2163_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2094_ __dut__._2094_/A1 __dut__._2094_/A2 __dut__._2093_/X VGND VGND VPWR
+ VPWR __dut__._2094_/X sky130_fd_sc_hd__a21o_4
XFILLER_80_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_38_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1947_ __dut__._2327_/A __dut__._2892_/Q VGND VGND VPWR VPWR __dut__._1947_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_140_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1878_ __dut__._1878_/A1 tie[166] __dut__._1877_/X VGND VGND VPWR VPWR __dut__._2858_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_106_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2289__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2285__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1921__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1752__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1504__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1280_ __dut__.__uuf__._1295_/A VGND VGND VPWR VPWR __dut__.__uuf__._1280_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2199__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1831__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2850_ clkbuf_5_6_0_tck/X __dut__._2850_/D __dut__._2402_/Y VGND VGND VPWR
+ VPWR __dut__._2850_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1616_ __dut__.__uuf__._1617_/A VGND VGND VPWR VPWR __dut__.__uuf__._1616_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1801_ __dut__._2213_/A __dut__._2819_/Q VGND VGND VPWR VPWR __dut__._1801_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1547_ __dut__.__uuf__._1558_/A VGND VGND VPWR VPWR __dut__.__uuf__._1547_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_107_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2781_ __dut__._2885_/CLK __dut__._2781_/D __dut__._2471_/Y VGND VGND VPWR
+ VPWR __dut__._2781_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1732_ __dut__._1910_/A1 tie[93] __dut__._1731_/X VGND VGND VPWR VPWR __dut__._2785_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1478_ __dut__.__uuf__._1478_/A VGND VGND VPWR VPWR __dut__.__uuf__._1478_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1663_ __dut__._1663_/A __dut__._2750_/Q VGND VGND VPWR VPWR __dut__._1663_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_131_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1594_ __dut__._1790_/A1 tie[24] __dut__._1593_/X VGND VGND VPWR VPWR __dut__._2716_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2215_ __dut__._2215_/A __dut__._2215_/B VGND VGND VPWR VPWR __dut__._2215_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2146_ __dut__._2146_/A1 __dut__._2146_/A2 __dut__._2145_/X VGND VGND VPWR
+ VPWR __dut__._2146_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_3_7_0_tck clkbuf_3_7_0_tck/A VGND VGND VPWR VPWR clkbuf_3_7_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2077_ __dut__._2213_/A __dut__._2077_/B VGND VGND VPWR VPWR __dut__._2077_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2572__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2695__CLK clkbuf_5_2_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_217_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2300__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2482__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_280 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1485_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_291 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2105_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1401_ __dut__.__uuf__._1401_/A VGND VGND VPWR VPWR __dut__.__uuf__._1401_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2381_ __dut__.__uuf__._2415_/CLK __dut__._2266_/X __dut__.__uuf__._1176_/X
+ VGND VGND VPWR VPWR __dut__._2267_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_117_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1332_ __dut__.__uuf__._1326_/X __dut__.__uuf__._1331_/X __dut__._2195_/B
+ __dut__.__uuf__._1326_/X VGND VGND VPWR VPWR __dut__._2194_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1263_ __dut__.__uuf__._1263_/A __dut__.__uuf__._1263_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1263_/Y sky130_fd_sc_hd__nand2_4
XFILLER_113_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1194_ __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR __dut__.__uuf__._1206_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_86_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2000_ __dut__._2000_/A1 __dut__._2000_/A2 __dut__._1999_/X VGND VGND VPWR
+ VPWR __dut__._2000_/X sky130_fd_sc_hd__a21o_4
XFILLER_42_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2392__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1716__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2833_ __dut__._2845_/CLK __dut__._2833_/D __dut__._2419_/Y VGND VGND VPWR
+ VPWR __dut__._2833_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2764_ __dut__._2865_/CLK __dut__._2764_/D __dut__._2488_/Y VGND VGND VPWR
+ VPWR __dut__._2764_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1715_ __dut__._1729_/A __dut__._2776_/Q VGND VGND VPWR VPWR __dut__._1715_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2695_ clkbuf_5_2_0_tck/X __dut__._2695_/D __dut__._2557_/Y VGND VGND VPWR
+ VPWR __dut__._2695_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1646_ __dut__._1646_/A1 tie[50] __dut__._1645_/X VGND VGND VPWR VPWR __dut__._2742_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1577_ __dut__._1793_/A __dut__._2707_/Q VGND VGND VPWR VPWR __dut__._1577_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1471__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2567__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2323__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0___dut__.__uuf__.__clk_source__/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2129_ __dut__._2149_/A __dut__._2129_/B VGND VGND VPWR VPWR __dut__._2129_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_146_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_167_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_334_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2477__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1950_ __dut__.__uuf__._1960_/A __dut__.__uuf__._1950_/B __dut__.__uuf__._1950_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1951_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1881_ __dut__._1308_/X VGND VGND VPWR VPWR __dut__.__uuf__._1885_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_32_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2860__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2364_ __dut__.__uuf__._2402_/CLK __dut__._2232_/X __dut__.__uuf__._1226_/X
+ VGND VGND VPWR VPWR __dut__._2233_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1315_ __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR __dut__.__uuf__._1315_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2295_ __dut__.__uuf__._2319_/CLK __dut__._2094_/X __dut__.__uuf__._1563_/X
+ VGND VGND VPWR VPWR __dut__._2095_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_143_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1500_ __dut__._1282_/Y mp[27] __dut__._1499_/X VGND VGND VPWR VPWR __dut__._1500_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._2480_ rst VGND VGND VPWR VPWR __dut__._2480_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1246_ __dut__.__uuf__._1341_/A VGND VGND VPWR VPWR __dut__.__uuf__._1429_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1431_ _234_/Y __dut__._2664_/Q VGND VGND VPWR VPWR __dut__._1431_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1177_ __dut__.__uuf__._1177_/A VGND VGND VPWR VPWR __dut__.__uuf__._1177_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1362_ __dut__._1362_/A1 __dut__._1360_/X __dut__._1361_/X VGND VGND VPWR
+ VPWR __dut__._2646_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1291__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2387__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1293_ __dut__._1293_/A __dut__._2628_/Q VGND VGND VPWR VPWR __dut__._1293_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_27_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_310_ _312_/CLK _310_/D trst VGND VGND VPWR VPWR _310_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_15_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_241_ _299_/Q _298_/Q _300_/Q VGND VGND VPWR VPWR _242_/D sky130_fd_sc_hd__or3_4
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_psn_inst_psn_buff_20_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_172_ _275_/Q _172_/B VGND VGND VPWR VPWR _274_/D sky130_fd_sc_hd__and2_4
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._2816_ clkbuf_5_0_0_tck/X __dut__._2816_/D __dut__._2436_/Y VGND VGND VPWR
+ VPWR __dut__._2816_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2747_ __dut__._2767_/CLK __dut__._2747_/D __dut__._2505_/Y VGND VGND VPWR
+ VPWR __dut__._2747_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2678_ __dut__._2680_/CLK __dut__._2678_/D __dut__._2574_/Y VGND VGND VPWR
+ VPWR __dut__._2678_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1629_ __dut__._1661_/A __dut__._2733_/Q VGND VGND VPWR VPWR __dut__._1629_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_92_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2297__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_284_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1100_ __dut__.__uuf__._1114_/A VGND VGND VPWR VPWR __dut__.__uuf__._1100_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2080_ VGND VGND VPWR VPWR __dut__.__uuf__._2080_/HI tie[25] sky130_fd_sc_hd__conb_1
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1031_ __dut__.__uuf__._2051_/A __dut__._1957_/B __dut__.__uuf__._1031_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1191_/A sky130_fd_sc_hd__or3_4
XFILLER_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1279__B2 __dut__.__uuf__._1040_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1933_ __dut__.__uuf__._1925_/A __dut__.__uuf__._1931_/B __dut__.__uuf__._1890_/X
+ VGND VGND VPWR VPWR __dut__._2038_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_52_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1864_ __dut__.__uuf__._1864_/A VGND VGND VPWR VPWR __dut__.__uuf__._1866_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1795_ __dut__._1991_/B __dut__._1997_/B VGND VGND VPWR VPWR __dut__.__uuf__._1796_/A
+ sky130_fd_sc_hd__and2_4
X__dut__._1980_ __dut__._1980_/A1 __dut__._1980_/A2 __dut__._1979_/X VGND VGND VPWR
+ VPWR __dut__._1980_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2416_ __dut__.__uuf__._2422_/CLK __dut__._2336_/X __dut__.__uuf__._1071_/X
+ VGND VGND VPWR VPWR __dut__._2337_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2344__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2347_ __dut__.__uuf__._2348_/CLK __dut__._2198_/X __dut__.__uuf__._1319_/X
+ VGND VGND VPWR VPWR __dut__._2199_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2601_ rst VGND VGND VPWR VPWR __dut__._2601_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2532_ rst VGND VGND VPWR VPWR __dut__._2532_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2278_ __dut__.__uuf__._2278_/CLK __dut__._2060_/X __dut__.__uuf__._1597_/X
+ VGND VGND VPWR VPWR __dut__._2061_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1229_ __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR __dut__.__uuf__._1229_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_87_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2463_ rst VGND VGND VPWR VPWR __dut__._2463_/Y sky130_fd_sc_hd__inv_2
X__dut__._2394_ rst VGND VGND VPWR VPWR __dut__._2394_/Y sky130_fd_sc_hd__inv_2
X__dut__._1414_ __dut__._1414_/A1 __dut__._1412_/X __dut__._1413_/X VGND VGND VPWR
+ VPWR __dut__._2659_/D sky130_fd_sc_hd__a21o_4
X__dut__._1345_ __dut__._1433_/A __dut__._2641_/Q VGND VGND VPWR VPWR __dut__._1345_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_224_ _298_/Q _224_/B VGND VGND VPWR VPWR _297_/D sky130_fd_sc_hd__and2_4
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_155_ _182_/A VGND VGND VPWR VPWR _163_/B sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2580__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1580_ __dut__.__uuf__._1564_/X __dut__.__uuf__._1890_/A __dut__._2087_/B
+ __dut__.__uuf__._1462_/A __dut__.__uuf__._1579_/X VGND VGND VPWR VPWR __dut__._2086_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_146_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2490__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2201_ VGND VGND VPWR VPWR __dut__.__uuf__._2201_/HI tie[146] sky130_fd_sc_hd__conb_1
XFILLER_142_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2132_ VGND VGND VPWR VPWR __dut__.__uuf__._2132_/HI tie[77] sky130_fd_sc_hd__conb_1
XFILLER_130_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2063_ VGND VGND VPWR VPWR __dut__.__uuf__._2063_/HI tie[8] sky130_fd_sc_hd__conb_1
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_109 psn_inst_psn_buff_99/A VGND VGND VPWR VPWR __dut__._1362_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_40_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1916_ __dut__._2035_/B __dut__._2041_/B __dut__.__uuf__._1915_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1917_/C sky130_fd_sc_hd__o21ai_4
XFILLER_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1847_ __dut__.__uuf__._1840_/A __dut__.__uuf__._1845_/B __dut__.__uuf__._1836_/X
+ VGND VGND VPWR VPWR __dut__._2006_/A2 sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._1368__A2 mc[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_24_0_tck clkbuf_5_25_0_tck/A VGND VGND VPWR VPWR _303_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1778_ __dut__.__uuf__._1778_/A VGND VGND VPWR VPWR __dut__.__uuf__._1780_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_125_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1963_ __dut__._2213_/A __dut__._1963_/B VGND VGND VPWR VPWR __dut__._1963_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_146_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1894_ __dut__._1894_/A1 prod[4] __dut__._1893_/X VGND VGND VPWR VPWR __dut__._2866_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_121_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1540__A2 mc[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2515_ rst VGND VGND VPWR VPWR __dut__._2515_/Y sky130_fd_sc_hd__inv_2
X__dut__._2446_ rst VGND VGND VPWR VPWR __dut__._2446_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2377_ rst VGND VGND VPWR VPWR __dut__._2377_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2575__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1328_ __dut__._1282_/Y mc[1] __dut__._1327_/X VGND VGND VPWR VPWR __dut__._1328_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_43_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_207_ _250_/Q _207_/B VGND VGND VPWR VPWR _207_/X sky130_fd_sc_hd__or2_4
XANTENNA___dut__._1919__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_138_ _236_/B _137_/B _137_/Y _127_/X VGND VGND VPWR VPWR _139_/A sky130_fd_sc_hd__a211o_4
XANTENNA___dut__._2308__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_247_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1286__A __dut__.__uuf__._1326_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2485__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1701_ __dut__._2343_/B __dut__.__uuf__._1695_/X __dut__._2279_/B
+ __dut__.__uuf__._1696_/X VGND VGND VPWR VPWR prod[24] sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1632_ __dut__.__uuf__._1636_/A VGND VGND VPWR VPWR __dut__.__uuf__._1632_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_119_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1829__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1563_ __dut__.__uuf__._1577_/A VGND VGND VPWR VPWR __dut__.__uuf__._1563_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_128_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1494_ __dut__.__uuf__._1494_/A VGND VGND VPWR VPWR __dut__.__uuf__._1494_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2115_ VGND VGND VPWR VPWR __dut__.__uuf__._2115_/HI tie[60] sky130_fd_sc_hd__conb_1
XFILLER_130_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2300_ __dut__._2356_/A1 __dut__._2300_/A2 __dut__._2299_/X VGND VGND VPWR
+ VPWR __dut__._2300_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1283__B _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2046_ __dut__.__uuf__._1742_/A __dut__.__uuf__._2044_/B __dut__.__uuf__._2044_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2047_/C sky130_fd_sc_hd__o21a_4
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2231_ __dut__._2313_/A __dut__._2231_/B VGND VGND VPWR VPWR __dut__._2231_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2395__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2162_ __dut__._2166_/A1 __dut__._2162_/A2 __dut__._2161_/X VGND VGND VPWR
+ VPWR __dut__._2162_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2093_ __dut__._2095_/A __dut__._2093_/B VGND VGND VPWR VPWR __dut__._2093_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_13_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1739__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1946_ __dut__._2328_/A1 prod[30] __dut__._1945_/X VGND VGND VPWR VPWR __dut__._2892_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_125_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1877_ __dut__._2213_/A __dut__._2857_/Q VGND VGND VPWR VPWR __dut__._1877_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_106_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2429_ rst VGND VGND VPWR VPWR __dut__._2429_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1504__A2 mc[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2817__CLK clkbuf_5_0_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1440__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1615_ __dut__.__uuf__._1617_/A VGND VGND VPWR VPWR __dut__.__uuf__._1615_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1546_ __dut__.__uuf__._1543_/X __dut__.__uuf__._1538_/X __dut__._2105_/B
+ __dut__.__uuf__._1527_/X __dut__.__uuf__._1545_/X VGND VGND VPWR VPWR __dut__._2104_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1800_ __dut__._1800_/A1 tie[127] __dut__._1799_/X VGND VGND VPWR VPWR __dut__._2819_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_107_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2780_ __dut__._2885_/CLK __dut__._2780_/D __dut__._2472_/Y VGND VGND VPWR
+ VPWR __dut__._2780_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1731_ __dut__._1733_/A __dut__._2784_/Q VGND VGND VPWR VPWR __dut__._1731_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1477_ __dut__.__uuf__._1494_/A VGND VGND VPWR VPWR __dut__.__uuf__._1477_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1662_ __dut__._1662_/A1 tie[58] __dut__._1661_/X VGND VGND VPWR VPWR __dut__._2750_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_103_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1593_ __dut__._1793_/A __dut__._2715_/Q VGND VGND VPWR VPWR __dut__._1593_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2029_ __dut__.__uuf__._2022_/A __dut__.__uuf__._2027_/B __dut__.__uuf__._1998_/X
+ VGND VGND VPWR VPWR __dut__._2074_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_45_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2214_ __dut__._2214_/A1 __dut__._2214_/A2 __dut__._2213_/X VGND VGND VPWR
+ VPWR __dut__._2214_/X sky130_fd_sc_hd__a21o_4
XFILLER_60_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2145_ __dut__._2149_/A __dut__._2145_/B VGND VGND VPWR VPWR __dut__._2145_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_50_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2076_ __dut__._2078_/A1 __dut__._2076_/A2 __dut__._2075_/X VGND VGND VPWR
+ VPWR __dut__._2076_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1929_ __dut__._2327_/A __dut__._2883_/Q VGND VGND VPWR VPWR __dut__._1929_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_136_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1564__A __dut__.__uuf__._1564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_112_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_281 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1481_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_270 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1661_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_292 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2103_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1379__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1400_ __dut__.__uuf__._1393_/X __dut__.__uuf__._1399_/X __dut__._2169_/B
+ __dut__.__uuf__._1393_/X VGND VGND VPWR VPWR __dut__._2168_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._2380_ __dut__.__uuf__._2412_/CLK __dut__._2264_/X __dut__.__uuf__._1180_/X
+ VGND VGND VPWR VPWR __dut__._2265_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_144_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1331_ __dut__.__uuf__._1330_/Y __dut__.__uuf__._1309_/X __dut__.__uuf__._1311_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1331_/X sky130_fd_sc_hd__o21a_4
XFILLER_116_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1262_ __dut__.__uuf__._1269_/A VGND VGND VPWR VPWR __dut__.__uuf__._1262_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1193_ __dut__.__uuf__._1192_/X __dut__.__uuf__._1188_/X __dut__._2257_/B
+ __dut__._2259_/B __dut__.__uuf__._1185_/X VGND VGND VPWR VPWR __dut__._2256_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_140_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2003__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2832_ __dut__._2845_/CLK __dut__._2832_/D __dut__._2420_/Y VGND VGND VPWR
+ VPWR __dut__._2832_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1529_ __dut__._1440_/X __dut__.__uuf__._1523_/X __dut__._2115_/B
+ __dut__.__uuf__._1528_/X VGND VGND VPWR VPWR __dut__.__uuf__._1529_/X sky130_fd_sc_hd__o22a_4
X__dut__._2763_ __dut__._2865_/CLK __dut__._2763_/D __dut__._2489_/Y VGND VGND VPWR
+ VPWR __dut__._2763_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1714_ __dut__._1726_/A1 tie[84] __dut__._1713_/X VGND VGND VPWR VPWR __dut__._2776_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._1649__A __dut__.__uuf__._1655_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2694_ clkbuf_5_2_0_tck/X __dut__._2694_/D __dut__._2558_/Y VGND VGND VPWR
+ VPWR __dut__._2694_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_psn_inst_psn_buff_98_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1645_ __dut__._1661_/A __dut__._2741_/Q VGND VGND VPWR VPWR __dut__._1645_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1576_ __dut__._1578_/A1 tie[15] __dut__._1575_/X VGND VGND VPWR VPWR __dut__._2707_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1404__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2583__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2128_ __dut__._2136_/A1 __dut__._2128_/A2 __dut__._2127_/X VGND VGND VPWR
+ VPWR __dut__._2128_/X sky130_fd_sc_hd__a21o_4
X__dut__._2059_ __dut__._2213_/A __dut__._2059_/B VGND VGND VPWR VPWR __dut__._2059_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1927__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_327_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1880_ __dut__.__uuf__._1988_/A VGND VGND VPWR VPWR __dut__.__uuf__._1931_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2298__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2493__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1946__A2 prod[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1837__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2363_ __dut__.__uuf__._2402_/CLK __dut__._2230_/X __dut__.__uuf__._1228_/X
+ VGND VGND VPWR VPWR __dut__._2231_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1314_ __dut__.__uuf__._1323_/A VGND VGND VPWR VPWR __dut__.__uuf__._1314_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_99_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0_tck clkbuf_3_7_0_tck/A VGND VGND VPWR VPWR clkbuf_3_6_0_tck/X sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._2294_ __dut__.__uuf__._2323_/CLK __dut__._2092_/X __dut__.__uuf__._1568_/X
+ VGND VGND VPWR VPWR __dut__._2093_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1245_ __dut__.__uuf__._1461_/A VGND VGND VPWR VPWR __dut__.__uuf__._1341_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_143_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1430_ __dut__._1430_/A1 __dut__._1428_/X __dut__._1429_/X VGND VGND VPWR
+ VPWR __dut__._2663_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1176_ __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR __dut__.__uuf__._1176_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1361_ __dut__._1361_/A __dut__._2645_/Q VGND VGND VPWR VPWR __dut__._1361_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_55_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1292_ __dut__._1282_/Y mc[11] __dut__._1291_/X VGND VGND VPWR VPWR __dut__._1292_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_240_ _240_/A VGND VGND VPWR VPWR _242_/C sky130_fd_sc_hd__inv_2
XFILLER_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_171_ _276_/Q _171_/B VGND VGND VPWR VPWR _275_/D sky130_fd_sc_hd__or2_4
XANTENNA_psn_inst_psn_buff_13_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1747__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2815_ clkbuf_5_0_0_tck/X __dut__._2815_/D __dut__._2437_/Y VGND VGND VPWR
+ VPWR __dut__._2815_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2746_ __dut__._2767_/CLK __dut__._2746_/D __dut__._2506_/Y VGND VGND VPWR
+ VPWR __dut__._2746_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2677_ __dut__._2680_/CLK __dut__._2677_/D __dut__._2575_/Y VGND VGND VPWR
+ VPWR __dut__._2677_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1628_ __dut__._1658_/A1 tie[41] __dut__._1627_/X VGND VGND VPWR VPWR __dut__._2733_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._2578__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1559_ __dut__._1611_/A __dut__._2698_/Q VGND VGND VPWR VPWR __dut__._1559_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_277_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2488__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1030_ __dut__.__uuf__._2051_/C VGND VGND VPWR VPWR __dut__.__uuf__._1031_/C
+ sky130_fd_sc_hd__inv_2
XFILLER_84_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__313__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1932_ __dut__.__uuf__._1932_/A VGND VGND VPWR VPWR __dut__._2040_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1863_ __dut__.__uuf__._1906_/A __dut__.__uuf__._1863_/B __dut__.__uuf__._1863_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1864_/A sky130_fd_sc_hd__or3_4
XFILLER_149_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1794_ __dut__._1536_/X VGND VGND VPWR VPWR __dut__.__uuf__._1798_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1451__A2 __dut__.__uuf__._1998_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2415_ __dut__.__uuf__._2415_/CLK __dut__._2334_/X __dut__.__uuf__._1075_/X
+ VGND VGND VPWR VPWR __dut__._2335_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._2313__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._2600_ rst VGND VGND VPWR VPWR __dut__._2600_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2346_ __dut__.__uuf__._2348_/CLK __dut__._2196_/X __dut__.__uuf__._1323_/X
+ VGND VGND VPWR VPWR __dut__._2197_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_120_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2531_ rst VGND VGND VPWR VPWR __dut__._2531_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2277_ __dut__.__uuf__._2278_/CLK __dut__._2058_/X __dut__.__uuf__._1598_/X
+ VGND VGND VPWR VPWR __dut__._2059_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2462_ rst VGND VGND VPWR VPWR __dut__._2462_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1228_ __dut__.__uuf__._1249_/A VGND VGND VPWR VPWR __dut__.__uuf__._1228_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2398__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1413_ __dut__._1433_/A __dut__._2658_/Q VGND VGND VPWR VPWR __dut__._1413_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2393_ rst VGND VGND VPWR VPWR __dut__._2393_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1159_ __dut__.__uuf__._1188_/A VGND VGND VPWR VPWR __dut__.__uuf__._1159_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1344_ __dut__._1282_/Y mc[23] __dut__._1343_/X VGND VGND VPWR VPWR __dut__._1344_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_103_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2280__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_223_ _299_/Q _297_/Q _231_/A VGND VGND VPWR VPWR _296_/D sky130_fd_sc_hd__o21a_4
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_154_ _192_/B VGND VGND VPWR VPWR _182_/A sky130_fd_sc_hd__inv_2
XFILLER_109_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2700__CLK clkbuf_5_2_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2729_ __dut__._2744_/CLK __dut__._2729_/D __dut__._2523_/Y VGND VGND VPWR
+ VPWR __dut__._2729_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1846__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2850__CLK clkbuf_5_6_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1387__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2200_ VGND VGND VPWR VPWR __dut__.__uuf__._2200_/HI tie[145] sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_1_0_0___dut__.__uuf__.__clk_source___A clkbuf_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2131_ VGND VGND VPWR VPWR __dut__.__uuf__._2131_/HI tie[76] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2062_ VGND VGND VPWR VPWR __dut__.__uuf__._2062_/HI tie[7] sky130_fd_sc_hd__conb_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2011__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1915_ __dut__.__uuf__._1915_/A VGND VGND VPWR VPWR __dut__.__uuf__._1915_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_25_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1846_ __dut__.__uuf__._1846_/A VGND VGND VPWR VPWR __dut__._2008_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_33_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1777_ __dut__.__uuf__._1798_/A __dut__.__uuf__._1777_/B __dut__.__uuf__._1777_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1778_/A sky130_fd_sc_hd__or3_4
XFILLER_137_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1962_ __dut__._1964_/A1 __dut__._1962_/A2 __dut__._1961_/X VGND VGND VPWR
+ VPWR __dut__._1962_/X sky130_fd_sc_hd__a21o_4
X__dut__._1893_ __dut__._2239_/A __dut__._2865_/Q VGND VGND VPWR VPWR __dut__._1893_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_133_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2329_ __dut__.__uuf__._2398_/CLK __dut__._2162_/X __dut__.__uuf__._1411_/X
+ VGND VGND VPWR VPWR __dut__._2163_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_58_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2514_ rst VGND VGND VPWR VPWR __dut__._2514_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1828__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_80_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2445_ rst VGND VGND VPWR VPWR __dut__._2445_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2376_ rst VGND VGND VPWR VPWR __dut__._2376_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1327_ _234_/Y __dut__._2638_/Q VGND VGND VPWR VPWR __dut__._1327_/X sky130_fd_sc_hd__and2_4
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2359__CLK __dut__.__uuf__._2402_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_43_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2591__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_206_ _210_/A VGND VGND VPWR VPWR _207_/B sky130_fd_sc_hd__inv_2
XFILLER_156_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_137_ _305_/Q _137_/B VGND VGND VPWR VPWR _137_/Y sky130_fd_sc_hd__nor2_4
XFILLER_99_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1935__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_142_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1700_ __dut__._2341_/B __dut__.__uuf__._1695_/X __dut__._2277_/B
+ __dut__.__uuf__._1696_/X VGND VGND VPWR VPWR prod[23] sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1631_ __dut__.__uuf__._1643_/A VGND VGND VPWR VPWR __dut__.__uuf__._1636_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_119_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1562_ __dut__.__uuf__._1581_/A VGND VGND VPWR VPWR __dut__.__uuf__._1577_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1493_ __dut__.__uuf__._1478_/X __dut__.__uuf__._1473_/X __dut__._2129_/B
+ __dut__.__uuf__._1484_/X __dut__.__uuf__._1492_/X VGND VGND VPWR VPWR __dut__._2128_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_115_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1845__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2114_ VGND VGND VPWR VPWR __dut__.__uuf__._2114_/HI tie[59] sky130_fd_sc_hd__conb_1
XFILLER_97_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2045_ __dut__.__uuf__._2045_/A VGND VGND VPWR VPWR __dut__.__uuf__._2047_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_151_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2230_ __dut__._2356_/A1 __dut__._2230_/A2 __dut__._2229_/X VGND VGND VPWR
+ VPWR __dut__._2230_/X sky130_fd_sc_hd__a21o_4
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2161_ __dut__._2167_/A __dut__._2161_/B VGND VGND VPWR VPWR __dut__._2161_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2092_ __dut__._2094_/A1 __dut__._2092_/A2 __dut__._2091_/X VGND VGND VPWR
+ VPWR __dut__._2092_/X sky130_fd_sc_hd__a21o_4
XFILLER_25_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1829_ __dut__.__uuf__._1829_/A VGND VGND VPWR VPWR __dut__.__uuf__._1829_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_40_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1945_ __dut__._2327_/A __dut__._2891_/Q VGND VGND VPWR VPWR __dut__._1945_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_118_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1876_ __dut__._1876_/A1 tie[165] __dut__._1875_/X VGND VGND VPWR VPWR __dut__._2857_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1755__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2428_ rst VGND VGND VPWR VPWR __dut__._2428_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2586__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2359_ rst VGND VGND VPWR VPWR __dut__._2359_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2496__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_5_23_0_tck clkbuf_5_23_0_tck/A VGND VGND VPWR VPWR _308_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1440__A2 mp[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1614_ __dut__.__uuf__._1617_/A VGND VGND VPWR VPWR __dut__.__uuf__._1614_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1545_ __dut__._1424_/X __dut__.__uuf__._1544_/X __dut__._2107_/B
+ __dut__.__uuf__._1528_/X VGND VGND VPWR VPWR __dut__.__uuf__._1545_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1730_ __dut__._1910_/A1 tie[92] __dut__._1729_/X VGND VGND VPWR VPWR __dut__._2784_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_104_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1575__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1476_ __dut__.__uuf__._1476_/A VGND VGND VPWR VPWR __dut__.__uuf__._1494_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_115_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1661_ __dut__._1661_/A __dut__._2749_/Q VGND VGND VPWR VPWR __dut__._1661_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1592_ __dut__._1790_/A1 tie[23] __dut__._1591_/X VGND VGND VPWR VPWR __dut__._2715_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2028_ __dut__.__uuf__._2028_/A VGND VGND VPWR VPWR __dut__._2076_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_57_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2213_ __dut__._2213_/A __dut__._2213_/B VGND VGND VPWR VPWR __dut__._2213_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_60_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2144_ __dut__._2144_/A1 __dut__._2144_/A2 __dut__._2143_/X VGND VGND VPWR
+ VPWR __dut__._2144_/X sky130_fd_sc_hd__a21o_4
XFILLER_111_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_43_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2075_ __dut__._2213_/A __dut__._2075_/B VGND VGND VPWR VPWR __dut__._2075_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_139_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1928_ __dut__._2328_/A1 prod[21] __dut__._1927_/X VGND VGND VPWR VPWR __dut__._2883_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1859_ __dut__._2213_/A __dut__._2848_/Q VGND VGND VPWR VPWR __dut__._1859_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_4_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_282 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1477_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_260 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1689_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_271 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1529_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA_psn_inst_psn_buff_105_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_293 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2101_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_145_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1330_ __dut__._2197_/B VGND VGND VPWR VPWR __dut__.__uuf__._1330_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_144_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1395__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1261_ __dut__.__uuf__._1259_/Y __dut__.__uuf__._1260_/X __dut__.__uuf__._1229_/X
+ __dut__._2223_/B __dut__.__uuf__._1247_/X VGND VGND VPWR VPWR __dut__._2222_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1192_ __dut__.__uuf__._1478_/A VGND VGND VPWR VPWR __dut__.__uuf__._1192_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_140_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._2831_ __dut__._2845_/CLK __dut__._2831_/D __dut__._2421_/Y VGND VGND VPWR
+ VPWR __dut__._2831_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2762_ __dut__._2865_/CLK __dut__._2762_/D __dut__._2490_/Y VGND VGND VPWR
+ VPWR __dut__._2762_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1528_ __dut__.__uuf__._1771_/A VGND VGND VPWR VPWR __dut__.__uuf__._1528_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1713_ __dut__._1729_/A __dut__._2775_/Q VGND VGND VPWR VPWR __dut__._1713_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2693_ clkbuf_5_2_0_tck/X __dut__._2693_/D __dut__._2559_/Y VGND VGND VPWR
+ VPWR __dut__._2693_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1459_ __dut__.__uuf__._1455_/X __dut__.__uuf__._1450_/X __dut__._2145_/B
+ __dut__.__uuf__._2050_/B __dut__.__uuf__._1458_/X VGND VGND VPWR VPWR __dut__._2144_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_89_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1644_ __dut__._1644_/A1 tie[49] __dut__._1643_/X VGND VGND VPWR VPWR __dut__._2741_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_103_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1575_ __dut__._1793_/A __dut__._2706_/Q VGND VGND VPWR VPWR __dut__._1575_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1404__A2 mp[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2127_ __dut__._2149_/A __dut__._2127_/B VGND VGND VPWR VPWR __dut__._2127_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2058_ __dut__._2058_/A1 __dut__._2058_/A2 __dut__._2057_/X VGND VGND VPWR
+ VPWR __dut__._2058_/X sky130_fd_sc_hd__a21o_4
XFILLER_41_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2807__CLK clkbuf_opt_1_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1340__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1943__A __dut__._2327_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2362_ __dut__.__uuf__._2402_/CLK __dut__._2228_/X __dut__.__uuf__._1231_/X
+ VGND VGND VPWR VPWR __dut__._2229_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_105_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2293_ __dut__.__uuf__._2323_/CLK __dut__._2090_/X __dut__.__uuf__._1571_/X
+ VGND VGND VPWR VPWR __dut__._2091_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1313_ __dut__.__uuf__._1298_/X __dut__.__uuf__._1312_/X __dut__._2203_/B
+ __dut__.__uuf__._1298_/X VGND VGND VPWR VPWR __dut__._2202_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1244_ __dut__.__uuf__._1244_/A __dut__.__uuf__._1307_/A VGND VGND
+ VPWR VPWR __dut__.__uuf__._1461_/A sky130_fd_sc_hd__or2_4
XANTENNA___dut__._1853__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1175_ __dut__.__uuf__._1162_/X __dut__.__uuf__._1174_/X __dut__._2269_/B
+ __dut__._2271_/B __dut__.__uuf__._1171_/X VGND VGND VPWR VPWR __dut__._2268_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_100_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1360_ __dut__._1282_/Y mc[27] __dut__._1359_/X VGND VGND VPWR VPWR __dut__._1360_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2242__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1291_ _234_/Y __dut__._2629_/Q VGND VGND VPWR VPWR __dut__._1291_/X sky130_fd_sc_hd__and2_4
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_tck_A tck VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_170_ _277_/Q _172_/B VGND VGND VPWR VPWR _276_/D sky130_fd_sc_hd__and2_4
XFILLER_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2814_ clkbuf_5_9_0_tck/X __dut__._2814_/D __dut__._2438_/Y VGND VGND VPWR
+ VPWR __dut__._2814_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2745_ __dut__._2767_/CLK __dut__._2745_/D __dut__._2507_/Y VGND VGND VPWR
+ VPWR __dut__._2745_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2676_ __dut__._2680_/CLK __dut__._2676_/D __dut__._2576_/Y VGND VGND VPWR
+ VPWR __dut__._2676_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1763__A __dut__._1853_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1627_ __dut__._1661_/A __dut__._2732_/Q VGND VGND VPWR VPWR __dut__._1627_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1558_ __dut__._1564_/A1 tie[6] __dut__._1557_/X VGND VGND VPWR VPWR __dut__._2698_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_73_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1489_ __dut__._1489_/A __dut__._2677_/Q VGND VGND VPWR VPWR __dut__._1489_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_93_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2594__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_299_ _312_/CLK _299_/D trst VGND VGND VPWR VPWR _299_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_172_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1931_ __dut__.__uuf__._1931_/A __dut__.__uuf__._1931_/B __dut__.__uuf__._1931_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1932_/A sky130_fd_sc_hd__or3_4
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1862_ __dut__._2015_/B __dut__._2021_/B __dut__.__uuf__._1861_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1863_/C sky130_fd_sc_hd__o21ai_4
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1793_ __dut__.__uuf__._1786_/A __dut__.__uuf__._1791_/B __dut__.__uuf__._1782_/X
+ VGND VGND VPWR VPWR __dut__._1986_/A2 sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._2009__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2414_ __dut__.__uuf__._2415_/CLK __dut__._2332_/X __dut__.__uuf__._1077_/X
+ VGND VGND VPWR VPWR __dut__._2333_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2345_ __dut__.__uuf__._2348_/CLK __dut__._2194_/X __dut__.__uuf__._1329_/X
+ VGND VGND VPWR VPWR __dut__._2195_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2530_ rst VGND VGND VPWR VPWR __dut__._2530_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2276_ __dut__.__uuf__._2278_/CLK __dut__._2056_/X __dut__.__uuf__._1599_/X
+ VGND VGND VPWR VPWR __dut__._2057_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_120_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2461_ rst VGND VGND VPWR VPWR __dut__._2461_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1304__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1227_ __dut__.__uuf__._1221_/X __dut__.__uuf__._1218_/X __dut__._2233_/B
+ __dut__._2235_/B __dut__.__uuf__._1215_/X VGND VGND VPWR VPWR __dut__._2232_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1412_ __dut__._1282_/Y mp[7] __dut__._1411_/X VGND VGND VPWR VPWR __dut__._1412_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1158_ __dut__.__uuf__._1161_/A VGND VGND VPWR VPWR __dut__.__uuf__._1158_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2392_ rst VGND VGND VPWR VPWR __dut__._2392_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1343_ _234_/Y __dut__._2642_/Q VGND VGND VPWR VPWR __dut__._1343_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1089_ __dut__.__uuf__._1089_/A VGND VGND VPWR VPWR __dut__.__uuf__._1655_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_103_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1662__B __dut__._1957_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_222_ _302_/Q _224_/B VGND VGND VPWR VPWR _295_/D sky130_fd_sc_hd__and2_4
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_153_ _236_/A _309_/Q _153_/C _240_/A VGND VGND VPWR VPWR _192_/B sky130_fd_sc_hd__or4_4
XFILLER_136_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2589__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2728_ __dut__._2744_/CLK __dut__._2728_/D __dut__._2524_/Y VGND VGND VPWR
+ VPWR __dut__._2728_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._2288__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_78_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2659_ __dut__._2661_/CLK __dut__._2659_/D __dut__._2593_/Y VGND VGND VPWR
+ VPWR __dut__._2659_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_tck clkbuf_3_5_0_tck/A VGND VGND VPWR VPWR clkbuf_3_5_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1782__A1 __dut__._2176_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2499__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2130_ VGND VGND VPWR VPWR __dut__.__uuf__._2130_/HI tie[75] sky130_fd_sc_hd__conb_1
XFILLER_124_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2061_ VGND VGND VPWR VPWR __dut__.__uuf__._2061_/HI tie[6] sky130_fd_sc_hd__conb_1
XFILLER_96_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1914_ __dut__._2035_/B __dut__._2041_/B VGND VGND VPWR VPWR __dut__.__uuf__._1915_/A
+ sky130_fd_sc_hd__and2_4
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1845_ __dut__.__uuf__._1877_/A __dut__.__uuf__._1845_/B __dut__.__uuf__._1845_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1846_/A sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1776_ __dut__._1983_/B __dut__._1989_/B __dut__.__uuf__._1775_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1777_/C sky130_fd_sc_hd__o21ai_4
XFILLER_137_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1961_ __dut__._2213_/A __dut__._1961_/B VGND VGND VPWR VPWR __dut__._1961_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_152_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1892_ __dut__._1892_/A1 prod[3] __dut__._1891_/X VGND VGND VPWR VPWR __dut__._2865_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_133_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2328_ __dut__.__uuf__._2398_/CLK __dut__._2160_/X __dut__.__uuf__._1417_/X
+ VGND VGND VPWR VPWR __dut__._2161_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_121_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2513_ rst VGND VGND VPWR VPWR __dut__._2513_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2259_ __dut__.__uuf__._2270_/CLK __dut__._2022_/X __dut__.__uuf__._1621_/X
+ VGND VGND VPWR VPWR __dut__._2023_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2444_ rst VGND VGND VPWR VPWR __dut__._2444_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2375_ rst VGND VGND VPWR VPWR __dut__._2375_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1326_ __dut__._1346_/A1 __dut__._1324_/X __dut__._1325_/X VGND VGND VPWR
+ VPWR __dut__._2637_/D sky130_fd_sc_hd__a21o_4
XFILLER_28_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1764__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_205_ _205_/A _248_/Q _247_/Q VGND VGND VPWR VPWR _210_/A sky130_fd_sc_hd__or3_4
XFILLER_156_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_136_ _309_/Q VGND VGND VPWR VPWR _236_/B sky130_fd_sc_hd__inv_2
XFILLER_7_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1516__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_135_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2303__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_302_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1630_ __dut__.__uuf__._1630_/A VGND VGND VPWR VPWR __dut__.__uuf__._1630_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1561_ __dut__.__uuf__._1543_/X __dut__.__uuf__._1559_/X __dut__._2097_/B
+ __dut__.__uuf__._1548_/X __dut__.__uuf__._1560_/X VGND VGND VPWR VPWR __dut__._2096_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_119_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1492_ __dut__._1476_/X __dut__.__uuf__._1480_/X __dut__._2131_/B
+ __dut__.__uuf__._1485_/X VGND VGND VPWR VPWR __dut__.__uuf__._1492_/X sky130_fd_sc_hd__o22a_4
XFILLER_115_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2113_ VGND VGND VPWR VPWR __dut__.__uuf__._2113_/HI tie[58] sky130_fd_sc_hd__conb_1
XFILLER_69_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2044_ __dut__.__uuf__._2044_/A __dut__.__uuf__._2044_/B __dut__.__uuf__._2044_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2045_/A sky130_fd_sc_hd__or3_4
XFILLER_151_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1861__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2160_ __dut__._2166_/A1 __dut__._2160_/A2 __dut__._2159_/X VGND VGND VPWR
+ VPWR __dut__._2160_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2091_ __dut__._2095_/A __dut__._2091_/B VGND VGND VPWR VPWR __dut__._2091_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1828_ __dut__._2003_/B __dut__._2009_/B VGND VGND VPWR VPWR __dut__.__uuf__._1829_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_40_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1746__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__264__CLK _270_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2840__CLK clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1759_ __dut__._1460_/X VGND VGND VPWR VPWR __dut__.__uuf__._1763_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_153_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1944_ __dut__._2338_/A1 prod[29] __dut__._1943_/X VGND VGND VPWR VPWR __dut__._2891_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_109_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1875_ __dut__._2213_/A __dut__._2856_/Q VGND VGND VPWR VPWR __dut__._1875_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_7_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1771__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2427_ rst VGND VGND VPWR VPWR __dut__._2427_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__232__A1 _304_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2358_ __dut__._1282_/Y clk __dut__._2357_/X VGND VGND VPWR VPWR __dut__._2358_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_16_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1309_ __dut__._1309_/A __dut__._2632_/Q VGND VGND VPWR VPWR __dut__._1309_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2289_ __dut__._2313_/A __dut__._2289_/B VGND VGND VPWR VPWR __dut__._2289_/X
+ sky130_fd_sc_hd__and2_4
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0___dut__.__uuf__.__clk_source__ clkbuf_4_9_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2372_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_144_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_252_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0___dut__.__uuf__.__clk_source__ clkbuf_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR clkbuf_2_1_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._2863__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1613_ __dut__.__uuf__._1617_/A VGND VGND VPWR VPWR __dut__.__uuf__._1613_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_135_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1544_ __dut__.__uuf__._1565_/A VGND VGND VPWR VPWR __dut__.__uuf__._1544_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1475_ __dut__.__uuf__._1455_/X __dut__.__uuf__._1473_/X __dut__._2137_/B
+ __dut__.__uuf__._1462_/X __dut__.__uuf__._1474_/X VGND VGND VPWR VPWR __dut__._2136_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_89_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1660_ __dut__._1660_/A1 tie[57] __dut__._1659_/X VGND VGND VPWR VPWR __dut__._2749_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1591_ __dut__._1793_/A __dut__._2714_/Q VGND VGND VPWR VPWR __dut__._1591_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2349__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1591__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2027_ __dut__.__uuf__._2037_/A __dut__.__uuf__._2027_/B __dut__.__uuf__._2027_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2028_/A sky130_fd_sc_hd__or3_4
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._2212_ __dut__._2214_/A1 __dut__._2212_/A2 __dut__._2211_/X VGND VGND VPWR
+ VPWR __dut__._2212_/X sky130_fd_sc_hd__a21o_4
X__dut__._2143_ __dut__._2149_/A __dut__._2143_/B VGND VGND VPWR VPWR __dut__._2143_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_111_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_36_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2074_ __dut__._2078_/A1 __dut__._2074_/A2 __dut__._2073_/X VGND VGND VPWR
+ VPWR __dut__._2074_/X sky130_fd_sc_hd__a21o_4
XFILLER_9_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1251__A1 __dut__.__uuf__._1229_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1927_ __dut__._2327_/A __dut__._2882_/Q VGND VGND VPWR VPWR __dut__._1927_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_107_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1858_ __dut__._1858_/A1 tie[156] __dut__._1857_/X VGND VGND VPWR VPWR __dut__._2848_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__290__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1789_ __dut__._1793_/A __dut__._2813_/Q VGND VGND VPWR VPWR __dut__._1789_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2597__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_250 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1901_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_261 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1687_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_272 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR psn_inst_psn_buff_325/A
+ sky130_fd_sc_hd__buf_8
XFILLER_31_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_294 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1361_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_283 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1473_/A
+ sky130_fd_sc_hd__buf_2
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__307__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1260_ __dut__._2223_/B __dut__.__uuf__._1260_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1260_/X sky130_fd_sc_hd__or2_4
X__dut__.__uuf__._1191_ __dut__.__uuf__._1191_/A VGND VGND VPWR VPWR __dut__.__uuf__._1478_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_140_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_3_0_tck_A clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._2830_ __dut__._2845_/CLK __dut__._2830_/D __dut__._2422_/Y VGND VGND VPWR
+ VPWR __dut__._2830_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2761_ __dut__._2865_/CLK __dut__._2761_/D __dut__._2491_/Y VGND VGND VPWR
+ VPWR __dut__._2761_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1527_ __dut__.__uuf__._1548_/A VGND VGND VPWR VPWR __dut__.__uuf__._1527_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2692_ clkbuf_5_2_0_tck/X __dut__._2692_/D __dut__._2560_/Y VGND VGND VPWR
+ VPWR __dut__._2692_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1712_ __dut__._1726_/A1 tie[83] __dut__._1711_/X VGND VGND VPWR VPWR __dut__._2775_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1458_ __dut__._1512_/X __dut__.__uuf__._1457_/X __dut__._2147_/B
+ __dut__.__uuf__._1438_/X VGND VGND VPWR VPWR __dut__.__uuf__._1458_/X sky130_fd_sc_hd__o22a_4
XFILLER_131_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1643_ __dut__._1643_/A __dut__._2740_/Q VGND VGND VPWR VPWR __dut__._1643_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1389_ __dut__.__uuf__._1414_/A VGND VGND VPWR VPWR __dut__.__uuf__._1389_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_106_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1574_ __dut__._1578_/A1 tie[14] __dut__._1573_/X VGND VGND VPWR VPWR __dut__._2706_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2126_ __dut__._2136_/A1 __dut__._2126_/A2 __dut__._2125_/X VGND VGND VPWR
+ VPWR __dut__._2126_/X sky130_fd_sc_hd__a21o_4
XFILLER_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2057_ __dut__._2213_/A __dut__._2057_/B VGND VGND VPWR VPWR __dut__._2057_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_5_22_0_tck clkbuf_5_23_0_tck/A VGND VGND VPWR VPWR __dut__._2892_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_142_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1340__A2 mc[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_215_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2356__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2361_ __dut__.__uuf__._2402_/CLK __dut__._2226_/X __dut__.__uuf__._1249_/X
+ VGND VGND VPWR VPWR __dut__._2227_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_145_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2292_ __dut__.__uuf__._2323_/CLK __dut__._2088_/X __dut__.__uuf__._1574_/X
+ VGND VGND VPWR VPWR __dut__._2089_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1312_ __dut__.__uuf__._1306_/Y __dut__.__uuf__._1309_/X __dut__.__uuf__._1311_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1312_/X sky130_fd_sc_hd__o21a_4
XFILLER_113_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1243_ __dut__.__uuf__._1456_/A VGND VGND VPWR VPWR __dut__.__uuf__._1307_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_99_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1766__A __dut__.__uuf__._2044_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1174_ __dut__.__uuf__._1188_/A VGND VGND VPWR VPWR __dut__.__uuf__._1174_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_39_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1290_ __dut__._1564_/A1 __dut__._1288_/X __dut__._1289_/X VGND VGND VPWR
+ VPWR __dut__._2628_/D sky130_fd_sc_hd__a21o_4
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2813_ clkbuf_5_9_0_tck/X __dut__._2813_/D __dut__._2439_/Y VGND VGND VPWR
+ VPWR __dut__._2813_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2205__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2744_ __dut__._2744_/CLK __dut__._2744_/D __dut__._2508_/Y VGND VGND VPWR
+ VPWR __dut__._2744_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._2675_ __dut__._2680_/CLK __dut__._2675_/D __dut__._2577_/Y VGND VGND VPWR
+ VPWR __dut__._2675_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1626_ __dut__._1626_/A1 tie[40] __dut__._1625_/X VGND VGND VPWR VPWR __dut__._2732_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_77_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1557_ __dut__._1611_/A __dut__._2697_/Q VGND VGND VPWR VPWR __dut__._1557_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_100_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1488_ __dut__._1282_/Y mp[24] __dut__._1487_/X VGND VGND VPWR VPWR __dut__._1488_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_93_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2109_ __dut__._2109_/A __dut__._2109_/B VGND VGND VPWR VPWR __dut__._2109_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_14_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_298_ _193_/A _298_/D trst VGND VGND VPWR VPWR _298_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2115__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_165_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_332_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1930_ __dut__.__uuf__._1929_/X __dut__.__uuf__._1927_/B __dut__.__uuf__._1927_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1931_/C sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1861_ __dut__.__uuf__._1861_/A VGND VGND VPWR VPWR __dut__.__uuf__._1861_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1792_ __dut__.__uuf__._1792_/A VGND VGND VPWR VPWR __dut__._1988_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_20_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2413_ __dut__.__uuf__._2415_/CLK __dut__._2330_/X __dut__.__uuf__._1079_/X
+ VGND VGND VPWR VPWR __dut__._2331_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2344_ __dut__.__uuf__._2348_/CLK __dut__._2192_/X __dut__.__uuf__._1333_/X
+ VGND VGND VPWR VPWR __dut__._2193_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_121_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2275_ __dut__.__uuf__._2278_/CLK __dut__._2054_/X __dut__.__uuf__._1601_/X
+ VGND VGND VPWR VPWR __dut__._2055_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2460_ rst VGND VGND VPWR VPWR __dut__._2460_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1304__A2 mc[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1226_ __dut__.__uuf__._1249_/A VGND VGND VPWR VPWR __dut__.__uuf__._1226_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1411_ _234_/Y __dut__._2659_/Q VGND VGND VPWR VPWR __dut__._1411_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1157_ __dut__.__uuf__._1147_/X __dut__.__uuf__._1144_/X __dut__._2281_/B
+ __dut__._2283_/B __dut__.__uuf__._1156_/X VGND VGND VPWR VPWR __dut__._2280_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_101_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_0_0_tck_A clkbuf_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2391_ rst VGND VGND VPWR VPWR __dut__._2391_/Y sky130_fd_sc_hd__inv_2
X__dut__._1342_ __dut__._1346_/A1 __dut__._1340_/X __dut__._1341_/X VGND VGND VPWR
+ VPWR __dut__._2641_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1088_ __dut__.__uuf__._1087_/X __dut__.__uuf__._1084_/X __dut__._2327_/B
+ __dut__._2329_/B __dut__.__uuf__._1081_/X VGND VGND VPWR VPWR __dut__._2326_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_55_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_221_ _229_/A _295_/Q VGND VGND VPWR VPWR _294_/D sky130_fd_sc_hd__and2_4
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_152_ _312_/Q _311_/Q VGND VGND VPWR VPWR _240_/A sky130_fd_sc_hd__or2_4
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2727_ __dut__._2744_/CLK __dut__._2727_/D __dut__._2525_/Y VGND VGND VPWR
+ VPWR __dut__._2727_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2658_ __dut__._2661_/CLK __dut__._2658_/D __dut__._2594_/Y VGND VGND VPWR
+ VPWR __dut__._2658_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1609_ __dut__._1793_/A __dut__._2723_/Q VGND VGND VPWR VPWR __dut__._1609_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_93_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2589_ rst VGND VGND VPWR VPWR __dut__._2589_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_1_0___dut__.__uuf__.__clk_source__ clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_3_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_119_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_282_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1534__A2 __dut__._1532_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2060_ VGND VGND VPWR VPWR __dut__.__uuf__._2060_/HI tie[5] sky130_fd_sc_hd__conb_1
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1913_ __dut__._1320_/X VGND VGND VPWR VPWR __dut__.__uuf__._1917_/B
+ sky130_fd_sc_hd__inv_2
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1844_ __dut__.__uuf__._1821_/X __dut__.__uuf__._1842_/B __dut__.__uuf__._1842_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1845_/C sky130_fd_sc_hd__o21a_4
XFILLER_40_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1859__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1775_ __dut__.__uuf__._1775_/A VGND VGND VPWR VPWR __dut__.__uuf__._1775_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1960_ __dut__._1960_/A1 __dut__._1960_/A2 __dut__._1959_/X VGND VGND VPWR
+ VPWR __dut__._1960_/X sky130_fd_sc_hd__a21o_4
XFILLER_137_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1891_ __dut__._2239_/A __dut__._2864_/Q VGND VGND VPWR VPWR __dut__._1891_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_133_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2327_ __dut__.__uuf__._2335_/CLK __dut__._2158_/X __dut__.__uuf__._1422_/X
+ VGND VGND VPWR VPWR __dut__._2159_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2512_ rst VGND VGND VPWR VPWR __dut__._2512_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2258_ __dut__.__uuf__._2278_/CLK __dut__._2020_/X __dut__.__uuf__._1622_/X
+ VGND VGND VPWR VPWR __dut__._2021_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_87_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1209_ __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR __dut__.__uuf__._1220_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._2443_ rst VGND VGND VPWR VPWR __dut__._2443_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2189_ VGND VGND VPWR VPWR __dut__.__uuf__._2189_/HI tie[134] sky130_fd_sc_hd__conb_1
X__dut__._2374_ rst VGND VGND VPWR VPWR __dut__._2374_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1325_ __dut__._1325_/A __dut__._2636_/Q VGND VGND VPWR VPWR __dut__._1325_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_28_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1769__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_204_ _246_/Q VGND VGND VPWR VPWR _205_/A sky130_fd_sc_hd__inv_2
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_135_ _310_/Q _137_/B _134_/X _127_/X VGND VGND VPWR VPWR _310_/D sky130_fd_sc_hd__a211o_4
XFILLER_152_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_15_0_tck clkbuf_3_7_0_tck/X VGND VGND VPWR VPWR clkbuf_5_31_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_99_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1516__A2 mp[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1951__B __dut__._2894_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_128_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1452__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1560_ __dut__._1404_/X __dut__.__uuf__._1544_/X __dut__._2099_/B
+ __dut__.__uuf__._1549_/X VGND VGND VPWR VPWR __dut__.__uuf__._1560_/X sky130_fd_sc_hd__o22a_4
XFILLER_119_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1491_ __dut__.__uuf__._1494_/A VGND VGND VPWR VPWR __dut__.__uuf__._1491_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2303__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2112_ VGND VGND VPWR VPWR __dut__.__uuf__._2112_/HI tie[57] sky130_fd_sc_hd__conb_1
XFILLER_69_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2043_ __dut__._2083_/B __dut__._1965_/B __dut__.__uuf__._2042_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._2044_/C sky130_fd_sc_hd__o21ai_4
XFILLER_57_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2090_ __dut__._2090_/A1 __dut__._2090_/A2 __dut__._2089_/X VGND VGND VPWR
+ VPWR __dut__._2090_/X sky130_fd_sc_hd__a21o_4
XFILLER_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1589__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1827_ __dut__._1288_/X VGND VGND VPWR VPWR __dut__.__uuf__._1831_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_138_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1758_ __dut__.__uuf__._1751_/A __dut__.__uuf__._1756_/B __dut__.__uuf__._1723_/X
+ VGND VGND VPWR VPWR __dut__._1974_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_21_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1943_ __dut__._2327_/A __dut__._2890_/Q VGND VGND VPWR VPWR __dut__._1943_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1689_ __dut__._1528_/X VGND VGND VPWR VPWR __dut__.__uuf__._1689_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1874_ __dut__._1874_/A1 tie[164] __dut__._1873_/X VGND VGND VPWR VPWR __dut__._2856_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_109_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2213__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_tck clkbuf_3_5_0_tck/A VGND VGND VPWR VPWR clkbuf_4_9_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_125_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2426_ rst VGND VGND VPWR VPWR __dut__._2426_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2357_ _234_/Y __dut__._2357_/B VGND VGND VPWR VPWR __dut__._2357_/X sky130_fd_sc_hd__and2_4
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1308_ __dut__._1282_/Y mc[15] __dut__._1307_/X VGND VGND VPWR VPWR __dut__._1308_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._2288_ __dut__._2356_/A1 __dut__._2288_/A2 __dut__._2287_/X VGND VGND VPWR
+ VPWR __dut__._2288_/X sky130_fd_sc_hd__a21o_4
XFILLER_71_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1499__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1859__A __dut__._1300_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2123__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1612_ __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR __dut__.__uuf__._1617_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_147_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1543_ __dut__.__uuf__._1564_/A VGND VGND VPWR VPWR __dut__.__uuf__._1543_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1474_ __dut__._1492_/X __dut__.__uuf__._1457_/X __dut__._2139_/B
+ __dut__.__uuf__._1463_/X VGND VGND VPWR VPWR __dut__.__uuf__._1474_/X sky130_fd_sc_hd__o22a_4
XFILLER_131_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1590_ __dut__._1790_/A1 tie[22] __dut__._1589_/X VGND VGND VPWR VPWR __dut__._2714_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_130_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2026_ __dut__.__uuf__._1983_/X __dut__.__uuf__._2024_/B __dut__.__uuf__._2024_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2027_/C sky130_fd_sc_hd__o21a_4
XFILLER_84_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2211_ __dut__._2213_/A __dut__._2211_/B VGND VGND VPWR VPWR __dut__._2211_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2142_ __dut__._2142_/A1 __dut__._2142_/A2 __dut__._2141_/X VGND VGND VPWR
+ VPWR __dut__._2142_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1416__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2073_ __dut__._2213_/A __dut__._2073_/B VGND VGND VPWR VPWR __dut__._2073_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_111_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_29_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1926_ __dut__._2328_/A1 prod[20] __dut__._1925_/X VGND VGND VPWR VPWR __dut__._2882_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_134_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1857_ __dut__._2213_/A __dut__._2847_/Q VGND VGND VPWR VPWR __dut__._1857_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_4_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1788_ __dut__._1790_/A1 tie[121] __dut__._1787_/X VGND VGND VPWR VPWR __dut__._2813_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2409_ rst VGND VGND VPWR VPWR __dut__._2409_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_240 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2259_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpsn_inst_psn_buff_251 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1899_/A
+ sky130_fd_sc_hd__buf_2
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_262 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1685_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_273 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1525_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_129_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_284 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1465_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_295 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2099_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_144_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1957__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_195_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1190_ __dut__.__uuf__._1190_/A VGND VGND VPWR VPWR __dut__.__uuf__._1190_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_112_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__254__CLK _308_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2830__CLK __dut__._2845_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1867__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1526_ __dut__.__uuf__._1537_/A VGND VGND VPWR VPWR __dut__.__uuf__._1526_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2316__CLK __dut__.__uuf__._2323_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_135_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2760_ __dut__._2865_/CLK __dut__._2760_/D __dut__._2492_/Y VGND VGND VPWR
+ VPWR __dut__._2760_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1711_ __dut__._1729_/A __dut__._2774_/Q VGND VGND VPWR VPWR __dut__._1711_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2691_ clkbuf_5_2_0_tck/X __dut__._2691_/D __dut__._2561_/Y VGND VGND VPWR
+ VPWR __dut__._2691_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1457_ __dut__.__uuf__._1578_/A VGND VGND VPWR VPWR __dut__.__uuf__._1457_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_104_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1642_ __dut__._1950_/A1 tie[48] __dut__._1641_/X VGND VGND VPWR VPWR __dut__._2740_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1388_ __dut__.__uuf__._1711_/A VGND VGND VPWR VPWR __dut__.__uuf__._1388_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_131_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1573_ __dut__._1793_/A __dut__._2705_/Q VGND VGND VPWR VPWR __dut__._1573_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_85_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2009_ __dut__.__uuf__._2002_/A __dut__.__uuf__._2007_/B __dut__.__uuf__._1998_/X
+ VGND VGND VPWR VPWR __dut__._2066_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_82_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2125_ __dut__._2149_/A __dut__._2125_/B VGND VGND VPWR VPWR __dut__._2125_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_26_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2056_ __dut__._2056_/A1 __dut__._2056_/A2 __dut__._2055_/X VGND VGND VPWR
+ VPWR __dut__._2056_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1777__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1909_ __dut__._2327_/A __dut__._2873_/Q VGND VGND VPWR VPWR __dut__._1909_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2889_ __dut__._2892_/CLK __dut__._2889_/D __dut__._2363_/Y VGND VGND VPWR
+ VPWR __dut__._2889_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2853__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2401__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_110_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2360_ __dut__.__uuf__._2402_/CLK __dut__._2224_/X __dut__.__uuf__._1254_/X
+ VGND VGND VPWR VPWR __dut__._2225_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_132_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2291_ __dut__.__uuf__._2355_/CLK __dut__._2086_/X __dut__.__uuf__._1577_/X
+ VGND VGND VPWR VPWR __dut__._2087_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1311_ __dut__.__uuf__._1337_/A VGND VGND VPWR VPWR __dut__.__uuf__._1311_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1242_ __dut__._2229_/B __dut__.__uuf__._1242_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1242_/X sky130_fd_sc_hd__or2_4
XFILLER_113_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2311__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1173_ __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR __dut__.__uuf__._1173_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_67_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2292__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1782__A __dut__.__uuf__._1890_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1597__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2812_ clkbuf_5_9_0_tck/X __dut__._2812_/D __dut__._2440_/Y VGND VGND VPWR
+ VPWR __dut__._2812_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2743_ __dut__._2744_/CLK __dut__._2743_/D __dut__._2509_/Y VGND VGND VPWR
+ VPWR __dut__._2743_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1509_ __dut__.__uuf__._1501_/X __dut__.__uuf__._1495_/X __dut__._2123_/B
+ __dut__.__uuf__._1506_/X __dut__.__uuf__._1508_/X VGND VGND VPWR VPWR __dut__._2122_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_117_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2674_ __dut__._2726_/CLK __dut__._2674_/D __dut__._2578_/Y VGND VGND VPWR
+ VPWR __dut__._2674_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1625_ __dut__._1661_/A __dut__._2731_/Q VGND VGND VPWR VPWR __dut__._1625_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_96_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1556_ __dut__._1564_/A1 tie[5] __dut__._1555_/X VGND VGND VPWR VPWR __dut__._2697_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_133_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1487_ _234_/Y __dut__._2678_/Q VGND VGND VPWR VPWR __dut__._1487_/X sky130_fd_sc_hd__and2_4
XFILLER_73_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2108_ __dut__._2108_/A1 __dut__._2108_/A2 __dut__._2107_/X VGND VGND VPWR
+ VPWR __dut__._2108_/X sky130_fd_sc_hd__a21o_4
XFILLER_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2039_ __dut__._2051_/A __dut__._2039_/B VGND VGND VPWR VPWR __dut__._2039_/X
+ sky130_fd_sc_hd__and2_4
X_297_ _312_/CLK _297_/D trst VGND VGND VPWR VPWR _297_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2131__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_158_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_325_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1860_ __dut__._2015_/B __dut__._2021_/B VGND VGND VPWR VPWR __dut__.__uuf__._1861_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1791_ __dut__.__uuf__._1823_/A __dut__.__uuf__._1791_/B __dut__.__uuf__._1791_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1792_/A sky130_fd_sc_hd__or3_4
XFILLER_149_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2412_ __dut__.__uuf__._2412_/CLK __dut__._2328_/X __dut__.__uuf__._1083_/X
+ VGND VGND VPWR VPWR __dut__._2329_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2343_ __dut__.__uuf__._2348_/CLK __dut__._2190_/X __dut__.__uuf__._1340_/X
+ VGND VGND VPWR VPWR __dut__._2191_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2274_ __dut__.__uuf__._2278_/CLK __dut__._2052_/X __dut__.__uuf__._1602_/X
+ VGND VGND VPWR VPWR __dut__._2053_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_87_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1225_ __dut__.__uuf__._1221_/X __dut__.__uuf__._1218_/X __dut__._2235_/B
+ __dut__._2237_/B __dut__.__uuf__._1215_/X VGND VGND VPWR VPWR __dut__._2234_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1410_ __dut__._1410_/A1 __dut__._1408_/X __dut__._1409_/X VGND VGND VPWR
+ VPWR __dut__._2658_/D sky130_fd_sc_hd__a21o_4
X__dut__._2390_ rst VGND VGND VPWR VPWR __dut__._2390_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1156_ __dut__.__uuf__._1215_/A VGND VGND VPWR VPWR __dut__.__uuf__._1156_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1341_ __dut__._1341_/A __dut__._2640_/Q VGND VGND VPWR VPWR __dut__._1341_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1087_ __dut__.__uuf__._1103_/A VGND VGND VPWR VPWR __dut__.__uuf__._1087_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_21_0_tck clkbuf_5_21_0_tck/A VGND VGND VPWR VPWR __dut__._2869_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_220_ _290_/Q _219_/A _217_/X VGND VGND VPWR VPWR _293_/D sky130_fd_sc_hd__o21a_4
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1989_ __dut__._1352_/X VGND VGND VPWR VPWR __dut__.__uuf__._1993_/B
+ sky130_fd_sc_hd__inv_2
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_151_ _300_/Q VGND VGND VPWR VPWR _153_/C sky130_fd_sc_hd__inv_2
XFILLER_7_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_11_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2861__D __dut__._2861_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2726_ __dut__._2726_/CLK __dut__._2726_/D __dut__._2526_/Y VGND VGND VPWR
+ VPWR __dut__._2726_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2657_ __dut__._2661_/CLK __dut__._2657_/D __dut__._2595_/Y VGND VGND VPWR
+ VPWR __dut__._2657_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1608_ __dut__._1610_/A1 tie[31] __dut__._1607_/X VGND VGND VPWR VPWR __dut__._2723_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2588_ rst VGND VGND VPWR VPWR __dut__._2588_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1539_ _234_/Y __dut__._2691_/Q VGND VGND VPWR VPWR __dut__._1539_/X sky130_fd_sc_hd__and2_4
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1965__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_275_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1912_ __dut__.__uuf__._1966_/A VGND VGND VPWR VPWR __dut__.__uuf__._1960_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_37_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1843_ __dut__.__uuf__._1843_/A VGND VGND VPWR VPWR __dut__.__uuf__._1845_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_33_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1774_ __dut__._1983_/B __dut__._1989_/B VGND VGND VPWR VPWR __dut__.__uuf__._1775_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_20_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1875__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1890_ __dut__._2238_/A1 prod[2] __dut__._1889_/X VGND VGND VPWR VPWR __dut__._2864_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_145_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2326_ __dut__.__uuf__._2335_/CLK __dut__._2156_/X __dut__.__uuf__._1426_/X
+ VGND VGND VPWR VPWR __dut__._2157_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._2511_ rst VGND VGND VPWR VPWR __dut__._2511_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2257_ __dut__.__uuf__._2270_/CLK __dut__._2018_/X __dut__.__uuf__._1623_/X
+ VGND VGND VPWR VPWR __dut__._2019_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_102_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1208_ __dut__.__uuf__._1207_/X __dut__.__uuf__._1204_/X __dut__._2247_/B
+ __dut__._2249_/B __dut__.__uuf__._1200_/X VGND VGND VPWR VPWR __dut__._2246_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._2442_ rst VGND VGND VPWR VPWR __dut__._2442_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2188_ VGND VGND VPWR VPWR __dut__.__uuf__._2188_/HI tie[133] sky130_fd_sc_hd__conb_1
XFILLER_75_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2373_ rst VGND VGND VPWR VPWR __dut__._2373_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1139_ __dut__.__uuf__._1133_/X __dut__.__uuf__._1130_/X __dut__._2293_/B
+ __dut__._2295_/B __dut__.__uuf__._1126_/X VGND VGND VPWR VPWR __dut__._2292_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_90_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1324_ __dut__._1282_/Y mc[19] __dut__._1323_/X VGND VGND VPWR VPWR __dut__._1324_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_59_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_203_ _244_/Q VGND VGND VPWR VPWR _203_/Y sky130_fd_sc_hd__inv_2
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_134_ _306_/Q _230_/A VGND VGND VPWR VPWR _134_/X sky130_fd_sc_hd__and2_4
XFILLER_137_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1785__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2709_ __dut__._2721_/CLK __dut__._2709_/D __dut__._2543_/Y VGND VGND VPWR
+ VPWR __dut__._2709_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1452__A2 mp[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1490_ __dut__.__uuf__._1478_/X __dut__.__uuf__._1473_/X __dut__._2131_/B
+ __dut__.__uuf__._1484_/X __dut__.__uuf__._1489_/X VGND VGND VPWR VPWR __dut__._2130_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_127_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2111_ VGND VGND VPWR VPWR __dut__.__uuf__._2111_/HI tie[56] sky130_fd_sc_hd__conb_1
X__dut__.__uuf__._2042_ __dut__.__uuf__._2042_/A VGND VGND VPWR VPWR __dut__.__uuf__._2042_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_111_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1826_ __dut__.__uuf__._1988_/A VGND VGND VPWR VPWR __dut__.__uuf__._1877_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1757_ __dut__.__uuf__._1757_/A VGND VGND VPWR VPWR __dut__._1976_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_153_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1942_ __dut__._2328_/A1 prod[28] __dut__._1941_/X VGND VGND VPWR VPWR __dut__._2890_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1688_ __dut__.__uuf__._1702_/A VGND VGND VPWR VPWR __dut__.__uuf__._1688_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1873_ __dut__._2213_/A __dut__._2855_/Q VGND VGND VPWR VPWR __dut__._1873_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_109_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2309_ __dut__.__uuf__._2323_/CLK __dut__._2122_/X __dut__.__uuf__._1505_/X
+ VGND VGND VPWR VPWR __dut__._2123_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2425_ rst VGND VGND VPWR VPWR __dut__._2425_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2356_ __dut__._2356_/A1 __dut__._2356_/A2 __dut__._2355_/X VGND VGND VPWR
+ VPWR __dut__._2356_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1307_ _234_/Y __dut__._2633_/Q VGND VGND VPWR VPWR __dut__._1307_/X sky130_fd_sc_hd__and2_4
X__dut__._2287_ __dut__._2313_/A __dut__._2287_/B VGND VGND VPWR VPWR __dut__._2287_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2404__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_140_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_238_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1611_ __dut__.__uuf__._1611_/A VGND VGND VPWR VPWR __dut__.__uuf__._1611_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1542_ __dut__.__uuf__._1558_/A VGND VGND VPWR VPWR __dut__.__uuf__._1542_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1473_ __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR __dut__.__uuf__._1473_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_116_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2025_ __dut__.__uuf__._2025_/A VGND VGND VPWR VPWR __dut__.__uuf__._2027_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._2210_ __dut__._2210_/A1 __dut__._2210_/A2 __dut__._2209_/X VGND VGND VPWR
+ VPWR __dut__._2210_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2245__CLK __dut__.__uuf__._2288_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_57_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2141_ __dut__._2149_/A __dut__._2141_/B VGND VGND VPWR VPWR __dut__._2141_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1416__A2 mc[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_14_0_tck clkbuf_3_7_0_tck/X VGND VGND VPWR VPWR clkbuf_5_29_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2072_ __dut__._2078_/A1 __dut__._2072_/A2 __dut__._2071_/X VGND VGND VPWR
+ VPWR __dut__._2072_/X sky130_fd_sc_hd__a21o_4
XFILLER_111_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1809_ __dut__.__uuf__._1852_/A __dut__.__uuf__._1809_/B __dut__.__uuf__._1809_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1810_/A sky130_fd_sc_hd__or3_4
XFILLER_154_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1925_ __dut__._2327_/A __dut__._2881_/Q VGND VGND VPWR VPWR __dut__._1925_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1856_ __dut__._1856_/A1 tie[155] __dut__._1855_/X VGND VGND VPWR VPWR __dut__._2847_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1352__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1787_ __dut__._1793_/A __dut__._2812_/Q VGND VGND VPWR VPWR __dut__._1787_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_122_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2408_ rst VGND VGND VPWR VPWR __dut__._2408_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0___dut__.__uuf__.__clk_source___A clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2339_ __dut__._2339_/A __dut__._2339_/B VGND VGND VPWR VPWR __dut__._2339_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1303__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_230 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2267_/A
+ sky130_fd_sc_hd__buf_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_241 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2257_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_263 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1673_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_252 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1897_/A
+ sky130_fd_sc_hd__buf_2
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_285 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1469_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_274 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1521_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_296 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._2097_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1957__B __dut__._1957_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_188_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1973__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1894__A2 prod[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._2309__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_tck clkbuf_3_3_0_tck/A VGND VGND VPWR VPWR clkbuf_4_7_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_136_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1525_ __dut__.__uuf__._1522_/X __dut__.__uuf__._1517_/X __dut__._2115_/B
+ __dut__.__uuf__._1506_/X __dut__.__uuf__._1524_/X VGND VGND VPWR VPWR __dut__._2114_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_135_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1710_ __dut__._1726_/A1 tie[82] __dut__._1709_/X VGND VGND VPWR VPWR __dut__._2774_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2690_ clkbuf_5_2_0_tck/X __dut__._2690_/D __dut__._2562_/Y VGND VGND VPWR
+ VPWR __dut__._2690_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1456_ __dut__.__uuf__._1456_/A VGND VGND VPWR VPWR __dut__.__uuf__._1578_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_150_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1883__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1387_ __dut__._2175_/B VGND VGND VPWR VPWR __dut__.__uuf__._1387_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1641_ __dut__._1641_/A __dut__._2739_/Q VGND VGND VPWR VPWR __dut__._1641_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_131_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1572_ __dut__._1572_/A1 tie[13] __dut__._1571_/X VGND VGND VPWR VPWR __dut__._2705_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_100_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2008_ __dut__.__uuf__._2008_/A VGND VGND VPWR VPWR __dut__._2068_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_122_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2124_ __dut__._2136_/A1 __dut__._2124_/A2 __dut__._2123_/X VGND VGND VPWR
+ VPWR __dut__._2124_/X sky130_fd_sc_hd__a21o_4
XFILLER_82_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_41_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2055_ __dut__._2213_/A __dut__._2055_/B VGND VGND VPWR VPWR __dut__._2055_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1908_ __dut__._1910_/A1 prod[11] __dut__._1907_/X VGND VGND VPWR VPWR __dut__._2873_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2888_ __dut__._2892_/CLK __dut__._2888_/D __dut__._2364_/Y VGND VGND VPWR
+ VPWR __dut__._2888_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1839_ __dut__._2213_/A __dut__._2838_/Q VGND VGND VPWR VPWR __dut__._1839_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_150_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1793__A __dut__._1793_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2129__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_103_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1310_ __dut__.__uuf__._1414_/A VGND VGND VPWR VPWR __dut__.__uuf__._1337_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2290_ __dut__.__uuf__._2355_/CLK __dut__._2084_/X __dut__.__uuf__._1582_/X
+ VGND VGND VPWR VPWR __dut__._2085_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_132_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1316__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1241_ __dut__.__uuf__._1241_/A __dut__.__uuf__._1241_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1241_/X sky130_fd_sc_hd__or2_4
XFILLER_113_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1172_ __dut__.__uuf__._1162_/X __dut__.__uuf__._1159_/X __dut__._2271_/B
+ __dut__._2273_/B __dut__.__uuf__._1171_/X VGND VGND VPWR VPWR __dut__._2270_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2811_ clkbuf_5_9_0_tck/X __dut__._2811_/D __dut__._2441_/Y VGND VGND VPWR
+ VPWR __dut__._2811_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2742_ __dut__._2894_/CLK __dut__._2742_/D __dut__._2510_/Y VGND VGND VPWR
+ VPWR __dut__._2742_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1508_ __dut__._1464_/X __dut__.__uuf__._1502_/X __dut__._2125_/B
+ __dut__.__uuf__._1507_/X VGND VGND VPWR VPWR __dut__.__uuf__._1508_/X sky130_fd_sc_hd__o22a_4
XFILLER_151_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1439_ __dut__.__uuf__._1437_/Y __dut__.__uuf__._1438_/X __dut__.__uuf__._1337_/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._1439_/X sky130_fd_sc_hd__o21a_4
XFILLER_132_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2673_ __dut__._2726_/CLK __dut__._2673_/D __dut__._2579_/Y VGND VGND VPWR
+ VPWR __dut__._2673_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2502__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1624_ __dut__._1624_/A1 tie[39] __dut__._1623_/X VGND VGND VPWR VPWR __dut__._2731_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1555_ __dut__._1555_/A __dut__._2696_/Q VGND VGND VPWR VPWR __dut__._1555_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_89_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1486_ __dut__._1486_/A1 __dut__._1484_/X __dut__._1485_/X VGND VGND VPWR
+ VPWR __dut__._2677_/D sky130_fd_sc_hd__a21o_4
XFILLER_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2107_ __dut__._2107_/A __dut__._2107_/B VGND VGND VPWR VPWR __dut__._2107_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._2038_ __dut__._2046_/A1 __dut__._2038_/A2 __dut__._2037_/X VGND VGND VPWR
+ VPWR __dut__._2038_/X sky130_fd_sc_hd__a21o_4
X_296_ _303_/CLK _296_/D trst VGND VGND VPWR VPWR _296_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_127_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2412__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2044__A __dut__.__uuf__._2044_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2306__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_52_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_220_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_318_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1790_ __dut__.__uuf__._1766_/X __dut__.__uuf__._1788_/B __dut__.__uuf__._1788_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1791_/C sky130_fd_sc_hd__o21a_4
XFILLER_149_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2411_ __dut__.__uuf__._2412_/CLK __dut__._2326_/X __dut__.__uuf__._1086_/X
+ VGND VGND VPWR VPWR __dut__._2327_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2342_ __dut__.__uuf__._2348_/CLK __dut__._2188_/X __dut__.__uuf__._1346_/X
+ VGND VGND VPWR VPWR __dut__._2189_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_133_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2273_ __dut__.__uuf__._2278_/CLK __dut__._2050_/X __dut__.__uuf__._1603_/X
+ VGND VGND VPWR VPWR __dut__._2051_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1224_ __dut__.__uuf__._1249_/A VGND VGND VPWR VPWR __dut__.__uuf__._1224_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_87_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1155_ __dut__.__uuf__._1244_/A VGND VGND VPWR VPWR __dut__.__uuf__._1215_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_101_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1340_ __dut__._1282_/Y mc[22] __dut__._1339_/X VGND VGND VPWR VPWR __dut__._1340_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1086_ __dut__.__uuf__._1086_/A VGND VGND VPWR VPWR __dut__.__uuf__._1086_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__267__CLK _271_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1988_ __dut__.__uuf__._1988_/A VGND VGND VPWR VPWR __dut__.__uuf__._2037_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2843__CLK clkbuf_opt_2_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_150_ _310_/Q VGND VGND VPWR VPWR _236_/A sky130_fd_sc_hd__inv_2
XFILLER_11_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1033__A __dut__.__uuf__._1564_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1528__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2725_ __dut__._2726_/CLK __dut__._2725_/D __dut__._2527_/Y VGND VGND VPWR
+ VPWR __dut__._2725_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2656_ __dut__._2661_/CLK __dut__._2656_/D __dut__._2596_/Y VGND VGND VPWR
+ VPWR __dut__._2656_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1607_ __dut__._1793_/A __dut__._2722_/Q VGND VGND VPWR VPWR __dut__._1607_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1700__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2587_ rst VGND VGND VPWR VPWR __dut__._2587_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1538_ __dut__._1538_/A1 __dut__._1536_/X __dut__._1537_/X VGND VGND VPWR
+ VPWR __dut__._2690_/D sky130_fd_sc_hd__a21o_4
XFILLER_73_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1469_ __dut__._1469_/A __dut__._2672_/Q VGND VGND VPWR VPWR __dut__._1469_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2407__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1311__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_279_ _288_/CLK _279_/D VGND VGND VPWR VPWR _279_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_155_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_170_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_268_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1981__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1911_ __dut__.__uuf__._1904_/A __dut__.__uuf__._1909_/B __dut__.__uuf__._1890_/X
+ VGND VGND VPWR VPWR __dut__._2030_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_25_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1118__A __dut__.__uuf__._1177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1842_ __dut__.__uuf__._1852_/A __dut__.__uuf__._1842_/B __dut__.__uuf__._1842_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1843_/A sky130_fd_sc_hd__or3_4
XANTENNA___dut__._1758__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1773_ __dut__._1504_/X VGND VGND VPWR VPWR __dut__.__uuf__._1777_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_138_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0___dut__.__uuf__.__clk_source__ clkbuf_2_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_133_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2325_ __dut__.__uuf__._2355_/CLK __dut__._2154_/X __dut__.__uuf__._1432_/X
+ VGND VGND VPWR VPWR __dut__._2155_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2510_ rst VGND VGND VPWR VPWR __dut__._2510_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2256_ __dut__.__uuf__._2278_/CLK __dut__._2016_/X __dut__.__uuf__._1624_/X
+ VGND VGND VPWR VPWR __dut__._2017_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2187_ VGND VGND VPWR VPWR __dut__.__uuf__._2187_/HI tie[132] sky130_fd_sc_hd__conb_1
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2441_ rst VGND VGND VPWR VPWR __dut__._2441_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1207_ __dut__.__uuf__._1478_/A VGND VGND VPWR VPWR __dut__.__uuf__._1207_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1138_ __dut__.__uuf__._1146_/A VGND VGND VPWR VPWR __dut__.__uuf__._1138_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_68_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2372_ rst VGND VGND VPWR VPWR __dut__._2372_/Y sky130_fd_sc_hd__inv_2
X__dut__._1323_ _234_/Y __dut__._2637_/Q VGND VGND VPWR VPWR __dut__._1323_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1069_ __dut__.__uuf__._1114_/A VGND VGND VPWR VPWR __dut__.__uuf__._1069_/X
+ sky130_fd_sc_hd__buf_2
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_202_ _202_/A VGND VGND VPWR VPWR _202_/X sky130_fd_sc_hd__buf_2
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_133_ _133_/A VGND VGND VPWR VPWR _311_/D sky130_fd_sc_hd__inv_2
XFILLER_137_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2174__A1 __dut__._2176_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2708_ __dut__._2721_/CLK __dut__._2708_/D __dut__._2544_/Y VGND VGND VPWR
+ VPWR __dut__._2708_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2639_ __dut__._2357_/B __dut__._2639_/D __dut__._2613_/Y VGND VGND VPWR
+ VPWR __dut__._2639_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2049__B1 __dut__.__uuf__._1038_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._2137__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_5_20_0_tck clkbuf_5_21_0_tck/A VGND VGND VPWR VPWR __dut__._2885_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2110_ VGND VGND VPWR VPWR __dut__.__uuf__._2110_/HI tie[55] sky130_fd_sc_hd__conb_1
XFILLER_130_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2041_ __dut__._2083_/B __dut__._1965_/B VGND VGND VPWR VPWR __dut__.__uuf__._2042_/A
+ sky130_fd_sc_hd__and2_4
XFILLER_111_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2600__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1825_ __dut__.__uuf__._1817_/A __dut__.__uuf__._1823_/B __dut__.__uuf__._1782_/X
+ VGND VGND VPWR VPWR __dut__._1998_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_100_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1756_ __dut__.__uuf__._1768_/A __dut__.__uuf__._1756_/B __dut__.__uuf__._1756_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1757_/A sky130_fd_sc_hd__or3_4
XFILLER_138_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1687_ __dut__._2323_/B __dut__.__uuf__._1681_/X __dut__._2259_/B
+ __dut__.__uuf__._1682_/X VGND VGND VPWR VPWR prod[14] sky130_fd_sc_hd__o22a_4
X__dut__._1941_ __dut__._2327_/A __dut__._2889_/Q VGND VGND VPWR VPWR __dut__._1941_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1872_ __dut__._1872_/A1 tie[163] __dut__._1871_/X VGND VGND VPWR VPWR __dut__._2855_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_119_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2308_ __dut__.__uuf__._2319_/CLK __dut__._2120_/X __dut__.__uuf__._1510_/X
+ VGND VGND VPWR VPWR __dut__._2121_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_125_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2239_ __dut__.__uuf__._2282_/CLK __dut__._1982_/X __dut__.__uuf__._1645_/X
+ VGND VGND VPWR VPWR __dut__._1983_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2510__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2424_ rst VGND VGND VPWR VPWR __dut__._2424_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2355_ __dut__._2355_/A __dut__._2355_/B VGND VGND VPWR VPWR __dut__._2355_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1306_ __dut__._1346_/A1 __dut__._1304_/X __dut__._1305_/X VGND VGND VPWR
+ VPWR __dut__._2632_/D sky130_fd_sc_hd__a21o_4
XFILLER_141_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2286_ __dut__._2356_/A1 __dut__._2286_/A2 __dut__._2285_/X VGND VGND VPWR
+ VPWR __dut__._2286_/X sky130_fd_sc_hd__a21o_4
XFILLER_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1221__A __dut__.__uuf__._1478_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2420__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_133_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_300_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1610_ __dut__.__uuf__._1611_/A VGND VGND VPWR VPWR __dut__.__uuf__._1610_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_147_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1541_ __dut__.__uuf__._1581_/A VGND VGND VPWR VPWR __dut__.__uuf__._1558_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_30_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1472_ __dut__.__uuf__._1472_/A VGND VGND VPWR VPWR __dut__.__uuf__._1472_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2310__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2024_ __dut__.__uuf__._2044_/A __dut__.__uuf__._2024_/B __dut__.__uuf__._2024_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2025_/A sky130_fd_sc_hd__or3_4
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2140_ __dut__._2140_/A1 __dut__._2140_/A2 __dut__._2139_/X VGND VGND VPWR
+ VPWR __dut__._2140_/X sky130_fd_sc_hd__a21o_4
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2071_ __dut__._2213_/A __dut__._2071_/B VGND VGND VPWR VPWR __dut__._2071_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_53_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1808_ __dut__._1995_/B __dut__._2001_/B __dut__.__uuf__._1807_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1809_/C sky130_fd_sc_hd__o21ai_4
XFILLER_139_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1739_ __dut__._1971_/B __dut__._1977_/B VGND VGND VPWR VPWR __dut__.__uuf__._1740_/A
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2505__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1924_ __dut__._2328_/A1 prod[19] __dut__._1923_/X VGND VGND VPWR VPWR __dut__._2881_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1855_ __dut__._2213_/A __dut__._2846_/Q VGND VGND VPWR VPWR __dut__._1855_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_134_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1352__A2 mc[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1786_ __dut__._1790_/A1 tie[120] __dut__._1785_/X VGND VGND VPWR VPWR __dut__._2812_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_96_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2407_ rst VGND VGND VPWR VPWR __dut__._2407_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_5_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2338_ __dut__._2338_/A1 __dut__._2338_/A2 __dut__._2337_/X VGND VGND VPWR
+ VPWR __dut__._2338_/X sky130_fd_sc_hd__a21o_4
X__dut__._2269_ __dut__._2269_/A __dut__._2269_/B VGND VGND VPWR VPWR __dut__._2269_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_32_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_231 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2317_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_220 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2271_/A
+ sky130_fd_sc_hd__buf_2
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_253 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2243_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_242 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2255_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_264 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1667_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_286 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1445_/A
+ sky130_fd_sc_hd__buf_2
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_275 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1517_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_297 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1365_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._2415__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_250_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1524_ __dut__._1444_/X __dut__.__uuf__._1523_/X __dut__._2117_/B
+ __dut__.__uuf__._1507_/X VGND VGND VPWR VPWR __dut__.__uuf__._1524_/X sky130_fd_sc_hd__o22a_4
XFILLER_151_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1455_ __dut__.__uuf__._1478_/A VGND VGND VPWR VPWR __dut__.__uuf__._1455_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1386_ __dut__.__uuf__._1401_/A VGND VGND VPWR VPWR __dut__.__uuf__._1386_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1640_ __dut__._1950_/A1 tie[47] __dut__._1639_/X VGND VGND VPWR VPWR __dut__._2739_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_131_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1571_ __dut__._1793_/A __dut__._2704_/Q VGND VGND VPWR VPWR __dut__._1571_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2007_ __dut__.__uuf__._2037_/A __dut__.__uuf__._2007_/B __dut__.__uuf__._2007_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2008_/A sky130_fd_sc_hd__or3_4
XFILLER_122_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2362__CLK __dut__.__uuf__._2402_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_73_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2123_ __dut__._2149_/A __dut__._2123_/B VGND VGND VPWR VPWR __dut__._2123_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_34_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._2054_ __dut__._2054_/A1 __dut__._2054_/A2 __dut__._2053_/X VGND VGND VPWR
+ VPWR __dut__._2054_/X sky130_fd_sc_hd__a21o_4
XFILLER_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2887_ __dut__._2892_/CLK __dut__._2887_/D __dut__._2365_/Y VGND VGND VPWR
+ VPWR __dut__._2887_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1907_ __dut__._1907_/A __dut__._2872_/Q VGND VGND VPWR VPWR __dut__._1907_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1838_ __dut__._2176_/A1 tie[146] __dut__._1837_/X VGND VGND VPWR VPWR __dut__._2838_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_122_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1769_ __dut__._2213_/A __dut__._2803_/Q VGND VGND VPWR VPWR __dut__._1769_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2145__A __dut__._2149_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2235__CLK __dut__.__uuf__._2282_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_298_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_4_0___dut__.__uuf__.__clk_source__ clkbuf_4_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2288_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_99_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_13_0_tck clkbuf_3_6_0_tck/X VGND VGND VPWR VPWR clkbuf_5_27_0_tck/A sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1316__A2 mc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1240_ __dut__.__uuf__._1242_/B VGND VGND VPWR VPWR __dut__.__uuf__._1241_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1171_ __dut__.__uuf__._1215_/A VGND VGND VPWR VPWR __dut__.__uuf__._1171_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_113_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._2810_ clkbuf_5_6_0_tck/X __dut__._2810_/D __dut__._2442_/Y VGND VGND VPWR
+ VPWR __dut__._2810_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._2055__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2741_ __dut__._2894_/CLK __dut__._2741_/D __dut__._2511_/Y VGND VGND VPWR
+ VPWR __dut__._2741_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1507_ __dut__.__uuf__._1507_/A VGND VGND VPWR VPWR __dut__.__uuf__._1507_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_104_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2672_ __dut__._2726_/CLK __dut__._2672_/D __dut__._2580_/Y VGND VGND VPWR
+ VPWR __dut__._2672_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1438_ __dut__.__uuf__._1507_/A VGND VGND VPWR VPWR __dut__.__uuf__._1438_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1623_ __dut__._1661_/A __dut__._2730_/Q VGND VGND VPWR VPWR __dut__._1623_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1369_ __dut__.__uuf__._1368_/Y __dut__.__uuf__._1362_/X __dut__.__uuf__._1363_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1369_/X sky130_fd_sc_hd__o21a_4
XFILLER_133_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1554_ __dut__._1554_/A1 tie[4] __dut__._1553_/X VGND VGND VPWR VPWR __dut__._2696_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_46_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1485_ __dut__._1485_/A __dut__._2676_/Q VGND VGND VPWR VPWR __dut__._1485_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_133_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2106_ __dut__._2106_/A1 __dut__._2106_/A2 __dut__._2105_/X VGND VGND VPWR
+ VPWR __dut__._2106_/X sky130_fd_sc_hd__a21o_4
X__dut__._2037_ __dut__._2051_/A __dut__._2037_/B VGND VGND VPWR VPWR __dut__._2037_/X
+ sky130_fd_sc_hd__and2_4
X_295_ _303_/CLK _295_/D trst VGND VGND VPWR VPWR _295_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_127_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_tck clkbuf_3_3_0_tck/A VGND VGND VPWR VPWR clkbuf_4_5_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1979__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_213_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2410_ __dut__.__uuf__._2412_/CLK __dut__._2324_/X __dut__.__uuf__._1092_/X
+ VGND VGND VPWR VPWR __dut__._2325_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_145_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2603__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2341_ __dut__.__uuf__._2348_/CLK __dut__._2186_/X __dut__.__uuf__._1350_/X
+ VGND VGND VPWR VPWR __dut__._2187_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2272_ __dut__.__uuf__._2278_/CLK __dut__._2048_/X __dut__.__uuf__._1604_/X
+ VGND VGND VPWR VPWR __dut__._2049_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_113_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2795__CLK _270_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1223_ __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR __dut__.__uuf__._1249_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_87_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1154_ __dut__.__uuf__._1161_/A VGND VGND VPWR VPWR __dut__.__uuf__._1154_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1085_ __dut__.__uuf__._1072_/X __dut__.__uuf__._1084_/X __dut__._2329_/B
+ __dut__._2331_/B __dut__.__uuf__._1081_/X VGND VGND VPWR VPWR __dut__._2328_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__300__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1889__A __dut__._2313_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2400__CLK __dut__.__uuf__._2402_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1987_ __dut__.__uuf__._1979_/A __dut__.__uuf__._1985_/B __dut__.__uuf__._1944_/X
+ VGND VGND VPWR VPWR __dut__._2058_/A2 sky130_fd_sc_hd__o21a_4
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1528__A2 prod_sel VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._2513__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2724_ clkbuf_5_8_0_tck/X __dut__._2724_/D __dut__._2528_/Y VGND VGND VPWR
+ VPWR __dut__._2724_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2655_ __dut__._2661_/CLK __dut__._2655_/D __dut__._2597_/Y VGND VGND VPWR
+ VPWR __dut__._2655_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1606_ __dut__._1610_/A1 tie[30] __dut__._1605_/X VGND VGND VPWR VPWR __dut__._2722_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2586_ rst VGND VGND VPWR VPWR __dut__._2586_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1537_ __dut__._1541_/A __dut__._2689_/Q VGND VGND VPWR VPWR __dut__._1537_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1464__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1468_ __dut__._1282_/Y mp[19] __dut__._1467_/X VGND VGND VPWR VPWR __dut__._1468_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_18_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1399_ _234_/Y __dut__._2656_/Q VGND VGND VPWR VPWR __dut__._1399_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1799__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_278_ _288_/CLK _278_/D VGND VGND VPWR VPWR _278_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2423__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_163_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_330_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1910_ __dut__.__uuf__._1910_/A VGND VGND VPWR VPWR __dut__._2032_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_25_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1841_ __dut__._2007_/B __dut__._2013_/B __dut__.__uuf__._1840_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._1842_/C sky130_fd_sc_hd__o21ai_4
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1772_ __dut__.__uuf__._1988_/A VGND VGND VPWR VPWR __dut__.__uuf__._1823_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_134_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2324_ __dut__.__uuf__._2355_/CLK __dut__._2152_/X __dut__.__uuf__._1436_/X
+ VGND VGND VPWR VPWR __dut__._2153_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1930__A2 prod[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2255_ __dut__.__uuf__._2278_/CLK __dut__._2014_/X __dut__.__uuf__._1626_/X
+ VGND VGND VPWR VPWR __dut__._2015_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_114_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2186_ VGND VGND VPWR VPWR __dut__.__uuf__._2186_/HI tie[131] sky130_fd_sc_hd__conb_1
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1206_ __dut__.__uuf__._1206_/A VGND VGND VPWR VPWR __dut__.__uuf__._1206_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._2440_ rst VGND VGND VPWR VPWR __dut__._2440_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1137_ __dut__.__uuf__._1133_/X __dut__.__uuf__._1130_/X __dut__._2295_/B
+ __dut__._2297_/B __dut__.__uuf__._1126_/X VGND VGND VPWR VPWR __dut__._2294_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_114_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2371_ rst VGND VGND VPWR VPWR __dut__._2371_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1322_ __dut__._1322_/A1 __dut__._1320_/X __dut__._1321_/X VGND VGND VPWR
+ VPWR __dut__._2636_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1068_ __dut__.__uuf__._1071_/A VGND VGND VPWR VPWR __dut__.__uuf__._1068_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_83_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2810__CLK clkbuf_5_6_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._2508__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_201_ _202_/A VGND VGND VPWR VPWR _201_/X sky130_fd_sc_hd__buf_2
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1044__A __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_132_ _130_/Y _230_/A _131_/Y _127_/X VGND VGND VPWR VPWR _133_/A sky130_fd_sc_hd__a211o_4
XFILLER_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2707_ clkbuf_5_0_0_tck/X __dut__._2707_/D __dut__._2545_/Y VGND VGND VPWR
+ VPWR __dut__._2707_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__293__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2638_ clkbuf_5_3_0_tck/X __dut__._2638_/D __dut__._2614_/Y VGND VGND VPWR
+ VPWR __dut__._2638_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2569_ rst VGND VGND VPWR VPWR __dut__._2569_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2418__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_280_A psn_inst_psn_buff_325/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2040_ __dut__._1376_/X VGND VGND VPWR VPWR __dut__.__uuf__._2044_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_111_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1676__A1 __dut__._1726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2833__CLK __dut__._2845_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1428__A1 __dut__._1282_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1129__A __dut__.__uuf__._1479_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1824_ __dut__.__uuf__._1824_/A VGND VGND VPWR VPWR __dut__._2000_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1755_ __dut__.__uuf__._1276_/X __dut__.__uuf__._1753_/B __dut__.__uuf__._1753_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1756_/C sky130_fd_sc_hd__o21a_4
XANTENNA___dut__.__uuf__._2319__CLK __dut__.__uuf__._2319_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1940_ __dut__._2328_/A1 prod[27] __dut__._1939_/X VGND VGND VPWR VPWR __dut__._2889_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1686_ __dut__._2321_/B __dut__.__uuf__._1681_/X __dut__._2257_/B
+ __dut__.__uuf__._1682_/X VGND VGND VPWR VPWR prod[13] sky130_fd_sc_hd__o22a_4
XFILLER_146_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1871_ __dut__._2213_/A __dut__._2854_/Q VGND VGND VPWR VPWR __dut__._1871_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_119_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2063__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2307_ __dut__.__uuf__._2319_/CLK __dut__._2118_/X __dut__.__uuf__._1513_/X
+ VGND VGND VPWR VPWR __dut__._2119_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2238_ __dut__.__uuf__._2282_/CLK __dut__._1980_/X __dut__.__uuf__._1646_/X
+ VGND VGND VPWR VPWR __dut__._1981_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_88_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2169_ VGND VGND VPWR VPWR __dut__.__uuf__._2169_/HI tie[114] sky130_fd_sc_hd__conb_1
XFILLER_125_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2423_ rst VGND VGND VPWR VPWR __dut__._2423_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1407__A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._2354_ __dut__._2356_/A1 __dut__._2354_/A2 __dut__._2353_/X VGND VGND VPWR
+ VPWR __dut__._2354_/X sky130_fd_sc_hd__a21o_4
XFILLER_141_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1305_ __dut__._1305_/A __dut__._2631_/Q VGND VGND VPWR VPWR __dut__._1305_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_64_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2285_ __dut__._2285_/A __dut__._2285_/B VGND VGND VPWR VPWR __dut__._2285_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2856__CLK clkbuf_5_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1830__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_126_A psn_inst_psn_buff_99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1987__A __dut__._2213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1540_ __dut__.__uuf__._1522_/X __dut__.__uuf__._1538_/X __dut__._2107_/B
+ __dut__.__uuf__._1527_/X __dut__.__uuf__._1539_/X VGND VGND VPWR VPWR __dut__._2106_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1471_ __dut__.__uuf__._1455_/X __dut__.__uuf__._1450_/X __dut__._2139_/B
+ __dut__.__uuf__._1462_/X __dut__.__uuf__._1470_/X VGND VGND VPWR VPWR __dut__._2138_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2611__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2023_ __dut__._2075_/B __dut__._2081_/B __dut__.__uuf__._2022_/Y
+ VGND VGND VPWR VPWR __dut__.__uuf__._2024_/C sky130_fd_sc_hd__o21ai_4
XFILLER_84_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2070_ __dut__._2070_/A1 __dut__._2070_/A2 __dut__._2069_/X VGND VGND VPWR
+ VPWR __dut__._2070_/X sky130_fd_sc_hd__a21o_4
XFILLER_80_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1807_ __dut__.__uuf__._1807_/A VGND VGND VPWR VPWR __dut__.__uuf__._1807_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_139_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1738_ __dut__._1372_/X VGND VGND VPWR VPWR __dut__.__uuf__._1742_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2291__CLK __dut__.__uuf__._2355_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_107_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1923_ __dut__._2327_/A __dut__._2880_/Q VGND VGND VPWR VPWR __dut__._1923_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1669_ __dut__._2295_/B __dut__.__uuf__._1666_/X __dut__._2231_/B
+ __dut__.__uuf__._1668_/X VGND VGND VPWR VPWR prod[0] sky130_fd_sc_hd__o22a_4
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1854_ __dut__._1854_/A1 tie[154] __dut__._1853_/X VGND VGND VPWR VPWR __dut__._2846_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_106_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1888__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._2521__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1785_ __dut__._1793_/A __dut__._2811_/Q VGND VGND VPWR VPWR __dut__._1785_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_121_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2406_ rst VGND VGND VPWR VPWR __dut__._2406_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2337_ __dut__._2337_/A __dut__._2337_/B VGND VGND VPWR VPWR __dut__._2337_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_45_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._2268_ __dut__._2268_/A1 __dut__._2268_/A2 __dut__._2267_/X VGND VGND VPWR
+ VPWR __dut__._2268_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1812__A1 __dut__._1854_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_210 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1817_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_221 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR psn_inst_psn_buff_228/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_254 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1709_/A
+ sky130_fd_sc_hd__buf_2
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_243 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR psn_inst_psn_buff_246/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_232 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._2319_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._2199_ __dut__._2213_/A __dut__._2199_/B VGND VGND VPWR VPWR __dut__._2199_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_276 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1513_/A
+ sky130_fd_sc_hd__buf_2
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_287 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1449_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_265 psn_inst_psn_buff_339/A VGND VGND VPWR VPWR __dut__._1665_/A
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_298 psn_inst_psn_buff_325/A VGND VGND VPWR VPWR __dut__._1417_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_129_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2431__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_243_A psn_inst_psn_buff_339/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2606__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1523_ __dut__.__uuf__._1565_/A VGND VGND VPWR VPWR __dut__.__uuf__._1523_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1454_ __dut__.__uuf__._1472_/A VGND VGND VPWR VPWR __dut__.__uuf__._1454_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1385_ __dut__.__uuf__._1378_/X __dut__.__uuf__._1384_/X __dut__._2175_/B
+ __dut__.__uuf__._1378_/X VGND VGND VPWR VPWR __dut__._2174_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1570_ __dut__._1570_/A1 tie[12] __dut__._1569_/X VGND VGND VPWR VPWR __dut__._2704_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_106_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2006_ __dut__.__uuf__._1983_/X __dut__.__uuf__._2004_/B __dut__.__uuf__._2004_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2007_/C sky130_fd_sc_hd__o21a_4
XFILLER_85_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2122_ __dut__._2136_/A1 __dut__._2122_/A2 __dut__._2121_/X VGND VGND VPWR
+ VPWR __dut__._2122_/X sky130_fd_sc_hd__a21o_4
XFILLER_81_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._2053_ __dut__._2213_/A __dut__._2053_/B VGND VGND VPWR VPWR __dut__._2053_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_41_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._2516__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_27_A __dut__._1772_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1906_ __dut__._1906_/A1 prod[10] __dut__._1905_/X VGND VGND VPWR VPWR __dut__._2872_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._2886_ __dut__._2892_/CLK __dut__._2886_/D __dut__._2366_/Y VGND VGND VPWR
+ VPWR __dut__._2886_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1837_ __dut__._1853_/A __dut__._2837_/Q VGND VGND VPWR VPWR __dut__._1837_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_135_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1768_ __dut__._1768_/A1 tie[111] __dut__._1767_/X VGND VGND VPWR VPWR __dut__._2803_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_110_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1699_ __dut__._1701_/A __dut__._2768_/Q VGND VGND VPWR VPWR __dut__._1699_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._2286__A1 __dut__._2356_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._2426__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_193_A psn_inst_psn_buff_193/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1170_ __dut__.__uuf__._1176_/A VGND VGND VPWR VPWR __dut__.__uuf__._1170_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_140_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

