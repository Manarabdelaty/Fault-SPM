VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spm_top
  CLASS BLOCK ;
  FOREIGN spm_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 297.880 300.000 298.480 ;
    END
  END done
  PIN mc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 0.720 300.000 1.320 ;
    END
  END mc[0]
  PIN mc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.160 300.000 23.760 ;
    END
  END mc[10]
  PIN mc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 25.880 300.000 26.480 ;
    END
  END mc[11]
  PIN mc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 27.920 300.000 28.520 ;
    END
  END mc[12]
  PIN mc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 30.640 300.000 31.240 ;
    END
  END mc[13]
  PIN mc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 32.680 300.000 33.280 ;
    END
  END mc[14]
  PIN mc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 34.720 300.000 35.320 ;
    END
  END mc[15]
  PIN mc[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 37.440 300.000 38.040 ;
    END
  END mc[16]
  PIN mc[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 39.480 300.000 40.080 ;
    END
  END mc[17]
  PIN mc[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 42.200 300.000 42.800 ;
    END
  END mc[18]
  PIN mc[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.240 300.000 44.840 ;
    END
  END mc[19]
  PIN mc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 2.760 300.000 3.360 ;
    END
  END mc[1]
  PIN mc[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 46.280 300.000 46.880 ;
    END
  END mc[20]
  PIN mc[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 49.000 300.000 49.600 ;
    END
  END mc[21]
  PIN mc[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 51.040 300.000 51.640 ;
    END
  END mc[22]
  PIN mc[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 53.760 300.000 54.360 ;
    END
  END mc[23]
  PIN mc[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 55.800 300.000 56.400 ;
    END
  END mc[24]
  PIN mc[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.840 300.000 58.440 ;
    END
  END mc[25]
  PIN mc[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 60.560 300.000 61.160 ;
    END
  END mc[26]
  PIN mc[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 62.600 300.000 63.200 ;
    END
  END mc[27]
  PIN mc[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 64.640 300.000 65.240 ;
    END
  END mc[28]
  PIN mc[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 67.360 300.000 67.960 ;
    END
  END mc[29]
  PIN mc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 4.800 300.000 5.400 ;
    END
  END mc[2]
  PIN mc[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 69.400 300.000 70.000 ;
    END
  END mc[30]
  PIN mc[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 72.120 300.000 72.720 ;
    END
  END mc[31]
  PIN mc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 7.520 300.000 8.120 ;
    END
  END mc[3]
  PIN mc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 9.560 300.000 10.160 ;
    END
  END mc[4]
  PIN mc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 11.600 300.000 12.200 ;
    END
  END mc[5]
  PIN mc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 14.320 300.000 14.920 ;
    END
  END mc[6]
  PIN mc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.360 300.000 16.960 ;
    END
  END mc[7]
  PIN mc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 19.080 300.000 19.680 ;
    END
  END mc[8]
  PIN mc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 21.120 300.000 21.720 ;
    END
  END mc[9]
  PIN mp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 74.160 300.000 74.760 ;
    END
  END mp[0]
  PIN mp[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 97.280 300.000 97.880 ;
    END
  END mp[10]
  PIN mp[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 99.320 300.000 99.920 ;
    END
  END mp[11]
  PIN mp[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 102.040 300.000 102.640 ;
    END
  END mp[12]
  PIN mp[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 104.080 300.000 104.680 ;
    END
  END mp[13]
  PIN mp[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 106.800 300.000 107.400 ;
    END
  END mp[14]
  PIN mp[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 108.840 300.000 109.440 ;
    END
  END mp[15]
  PIN mp[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 110.880 300.000 111.480 ;
    END
  END mp[16]
  PIN mp[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 113.600 300.000 114.200 ;
    END
  END mp[17]
  PIN mp[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 115.640 300.000 116.240 ;
    END
  END mp[18]
  PIN mp[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 118.360 300.000 118.960 ;
    END
  END mp[19]
  PIN mp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.200 300.000 76.800 ;
    END
  END mp[1]
  PIN mp[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 120.400 300.000 121.000 ;
    END
  END mp[20]
  PIN mp[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.440 300.000 123.040 ;
    END
  END mp[21]
  PIN mp[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.160 300.000 125.760 ;
    END
  END mp[22]
  PIN mp[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 127.200 300.000 127.800 ;
    END
  END mp[23]
  PIN mp[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 129.240 300.000 129.840 ;
    END
  END mp[24]
  PIN mp[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 131.960 300.000 132.560 ;
    END
  END mp[25]
  PIN mp[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 134.000 300.000 134.600 ;
    END
  END mp[26]
  PIN mp[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.720 300.000 137.320 ;
    END
  END mp[27]
  PIN mp[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 138.760 300.000 139.360 ;
    END
  END mp[28]
  PIN mp[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 140.800 300.000 141.400 ;
    END
  END mp[29]
  PIN mp[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 78.920 300.000 79.520 ;
    END
  END mp[2]
  PIN mp[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 143.520 300.000 144.120 ;
    END
  END mp[30]
  PIN mp[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 145.560 300.000 146.160 ;
    END
  END mp[31]
  PIN mp[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 80.960 300.000 81.560 ;
    END
  END mp[3]
  PIN mp[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 83.680 300.000 84.280 ;
    END
  END mp[4]
  PIN mp[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 85.720 300.000 86.320 ;
    END
  END mp[5]
  PIN mp[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 87.760 300.000 88.360 ;
    END
  END mp[6]
  PIN mp[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 90.480 300.000 91.080 ;
    END
  END mp[7]
  PIN mp[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 92.520 300.000 93.120 ;
    END
  END mp[8]
  PIN mp[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 95.240 300.000 95.840 ;
    END
  END mp[9]
  PIN prod[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.280 300.000 148.880 ;
    END
  END prod[0]
  PIN prod[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 171.400 300.000 172.000 ;
    END
  END prod[10]
  PIN prod[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 173.440 300.000 174.040 ;
    END
  END prod[11]
  PIN prod[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 175.480 300.000 176.080 ;
    END
  END prod[12]
  PIN prod[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 178.200 300.000 178.800 ;
    END
  END prod[13]
  PIN prod[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 180.240 300.000 180.840 ;
    END
  END prod[14]
  PIN prod[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.280 300.000 182.880 ;
    END
  END prod[15]
  PIN prod[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 185.000 300.000 185.600 ;
    END
  END prod[16]
  PIN prod[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 187.040 300.000 187.640 ;
    END
  END prod[17]
  PIN prod[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 189.760 300.000 190.360 ;
    END
  END prod[18]
  PIN prod[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 191.800 300.000 192.400 ;
    END
  END prod[19]
  PIN prod[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 150.320 300.000 150.920 ;
    END
  END prod[1]
  PIN prod[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 193.840 300.000 194.440 ;
    END
  END prod[20]
  PIN prod[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 196.560 300.000 197.160 ;
    END
  END prod[21]
  PIN prod[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 198.600 300.000 199.200 ;
    END
  END prod[22]
  PIN prod[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.320 300.000 201.920 ;
    END
  END prod[23]
  PIN prod[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 203.360 300.000 203.960 ;
    END
  END prod[24]
  PIN prod[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.400 300.000 206.000 ;
    END
  END prod[25]
  PIN prod[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 208.120 300.000 208.720 ;
    END
  END prod[26]
  PIN prod[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 210.160 300.000 210.760 ;
    END
  END prod[27]
  PIN prod[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 212.880 300.000 213.480 ;
    END
  END prod[28]
  PIN prod[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 214.920 300.000 215.520 ;
    END
  END prod[29]
  PIN prod[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 152.360 300.000 152.960 ;
    END
  END prod[2]
  PIN prod[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 216.960 300.000 217.560 ;
    END
  END prod[30]
  PIN prod[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 219.680 300.000 220.280 ;
    END
  END prod[31]
  PIN prod[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.720 300.000 222.320 ;
    END
  END prod[32]
  PIN prod[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.440 300.000 225.040 ;
    END
  END prod[33]
  PIN prod[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 226.480 300.000 227.080 ;
    END
  END prod[34]
  PIN prod[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 228.520 300.000 229.120 ;
    END
  END prod[35]
  PIN prod[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 231.240 300.000 231.840 ;
    END
  END prod[36]
  PIN prod[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 233.280 300.000 233.880 ;
    END
  END prod[37]
  PIN prod[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 236.000 300.000 236.600 ;
    END
  END prod[38]
  PIN prod[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 238.040 300.000 238.640 ;
    END
  END prod[39]
  PIN prod[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 155.080 300.000 155.680 ;
    END
  END prod[3]
  PIN prod[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 240.080 300.000 240.680 ;
    END
  END prod[40]
  PIN prod[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 242.800 300.000 243.400 ;
    END
  END prod[41]
  PIN prod[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.840 300.000 245.440 ;
    END
  END prod[42]
  PIN prod[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 246.880 300.000 247.480 ;
    END
  END prod[43]
  PIN prod[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 249.600 300.000 250.200 ;
    END
  END prod[44]
  PIN prod[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 251.640 300.000 252.240 ;
    END
  END prod[45]
  PIN prod[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 254.360 300.000 254.960 ;
    END
  END prod[46]
  PIN prod[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 256.400 300.000 257.000 ;
    END
  END prod[47]
  PIN prod[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.440 300.000 259.040 ;
    END
  END prod[48]
  PIN prod[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 261.160 300.000 261.760 ;
    END
  END prod[49]
  PIN prod[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 157.120 300.000 157.720 ;
    END
  END prod[4]
  PIN prod[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 263.200 300.000 263.800 ;
    END
  END prod[50]
  PIN prod[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 265.920 300.000 266.520 ;
    END
  END prod[51]
  PIN prod[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 267.960 300.000 268.560 ;
    END
  END prod[52]
  PIN prod[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 270.000 300.000 270.600 ;
    END
  END prod[53]
  PIN prod[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 272.720 300.000 273.320 ;
    END
  END prod[54]
  PIN prod[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 274.760 300.000 275.360 ;
    END
  END prod[55]
  PIN prod[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.480 300.000 278.080 ;
    END
  END prod[56]
  PIN prod[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 279.520 300.000 280.120 ;
    END
  END prod[57]
  PIN prod[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 281.560 300.000 282.160 ;
    END
  END prod[58]
  PIN prod[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 284.280 300.000 284.880 ;
    END
  END prod[59]
  PIN prod[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 159.840 300.000 160.440 ;
    END
  END prod[5]
  PIN prod[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 286.320 300.000 286.920 ;
    END
  END prod[60]
  PIN prod[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.040 300.000 289.640 ;
    END
  END prod[61]
  PIN prod[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 291.080 300.000 291.680 ;
    END
  END prod[62]
  PIN prod[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 293.120 300.000 293.720 ;
    END
  END prod[63]
  PIN prod[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 161.880 300.000 162.480 ;
    END
  END prod[6]
  PIN prod[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 163.920 300.000 164.520 ;
    END
  END prod[7]
  PIN prod[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 166.640 300.000 167.240 ;
    END
  END prod[8]
  PIN prod[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 168.680 300.000 169.280 ;
    END
  END prod[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END rst
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 295.840 300.000 296.440 ;
    END
  END start
  PIN tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END tck
  PIN tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END tdi
  PIN tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END tdo
  PIN tdo_paden_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END tdo_paden_o
  PIN tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END tms
  PIN trst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 296.000 150.330 300.000 ;
    END
  END trst
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 295.175 288.405 ;
      LAYER met1 ;
        RECT 5.520 9.560 295.250 288.560 ;
      LAYER met2 ;
        RECT 15.270 295.720 149.770 298.365 ;
        RECT 150.610 295.720 295.230 298.365 ;
        RECT 15.270 4.280 295.230 295.720 ;
        RECT 15.270 0.835 29.710 4.280 ;
        RECT 30.550 0.835 89.510 4.280 ;
        RECT 90.350 0.835 149.310 4.280 ;
        RECT 150.150 0.835 209.570 4.280 ;
        RECT 210.410 0.835 269.370 4.280 ;
        RECT 270.210 0.835 295.230 4.280 ;
      LAYER met3 ;
        RECT 4.000 297.480 295.600 298.345 ;
        RECT 4.000 296.840 296.000 297.480 ;
        RECT 4.000 295.440 295.600 296.840 ;
        RECT 4.000 294.120 296.000 295.440 ;
        RECT 4.000 292.720 295.600 294.120 ;
        RECT 4.000 292.080 296.000 292.720 ;
        RECT 4.000 290.680 295.600 292.080 ;
        RECT 4.000 290.040 296.000 290.680 ;
        RECT 4.000 288.640 295.600 290.040 ;
        RECT 4.000 287.320 296.000 288.640 ;
        RECT 4.000 285.920 295.600 287.320 ;
        RECT 4.000 285.280 296.000 285.920 ;
        RECT 4.000 283.880 295.600 285.280 ;
        RECT 4.000 282.560 296.000 283.880 ;
        RECT 4.000 281.160 295.600 282.560 ;
        RECT 4.000 280.520 296.000 281.160 ;
        RECT 4.000 279.120 295.600 280.520 ;
        RECT 4.000 278.480 296.000 279.120 ;
        RECT 4.000 277.080 295.600 278.480 ;
        RECT 4.000 275.760 296.000 277.080 ;
        RECT 4.000 274.360 295.600 275.760 ;
        RECT 4.000 273.720 296.000 274.360 ;
        RECT 4.000 272.320 295.600 273.720 ;
        RECT 4.000 271.000 296.000 272.320 ;
        RECT 4.000 269.600 295.600 271.000 ;
        RECT 4.000 268.960 296.000 269.600 ;
        RECT 4.000 267.560 295.600 268.960 ;
        RECT 4.000 266.920 296.000 267.560 ;
        RECT 4.000 265.520 295.600 266.920 ;
        RECT 4.000 264.200 296.000 265.520 ;
        RECT 4.000 262.800 295.600 264.200 ;
        RECT 4.000 262.160 296.000 262.800 ;
        RECT 4.000 260.760 295.600 262.160 ;
        RECT 4.000 259.440 296.000 260.760 ;
        RECT 4.000 258.040 295.600 259.440 ;
        RECT 4.000 257.400 296.000 258.040 ;
        RECT 4.000 256.000 295.600 257.400 ;
        RECT 4.000 255.360 296.000 256.000 ;
        RECT 4.000 253.960 295.600 255.360 ;
        RECT 4.000 252.640 296.000 253.960 ;
        RECT 4.000 251.240 295.600 252.640 ;
        RECT 4.000 250.600 296.000 251.240 ;
        RECT 4.000 249.200 295.600 250.600 ;
        RECT 4.000 247.880 296.000 249.200 ;
        RECT 4.000 246.480 295.600 247.880 ;
        RECT 4.000 245.840 296.000 246.480 ;
        RECT 4.000 244.440 295.600 245.840 ;
        RECT 4.000 243.800 296.000 244.440 ;
        RECT 4.000 242.400 295.600 243.800 ;
        RECT 4.000 241.080 296.000 242.400 ;
        RECT 4.000 239.680 295.600 241.080 ;
        RECT 4.000 239.040 296.000 239.680 ;
        RECT 4.000 237.640 295.600 239.040 ;
        RECT 4.000 237.000 296.000 237.640 ;
        RECT 4.000 235.600 295.600 237.000 ;
        RECT 4.000 234.280 296.000 235.600 ;
        RECT 4.000 232.880 295.600 234.280 ;
        RECT 4.000 232.240 296.000 232.880 ;
        RECT 4.000 230.840 295.600 232.240 ;
        RECT 4.000 229.520 296.000 230.840 ;
        RECT 4.000 228.120 295.600 229.520 ;
        RECT 4.000 227.480 296.000 228.120 ;
        RECT 4.000 226.080 295.600 227.480 ;
        RECT 4.000 225.440 296.000 226.080 ;
        RECT 4.400 224.040 295.600 225.440 ;
        RECT 4.000 222.720 296.000 224.040 ;
        RECT 4.000 221.320 295.600 222.720 ;
        RECT 4.000 220.680 296.000 221.320 ;
        RECT 4.000 219.280 295.600 220.680 ;
        RECT 4.000 217.960 296.000 219.280 ;
        RECT 4.000 216.560 295.600 217.960 ;
        RECT 4.000 215.920 296.000 216.560 ;
        RECT 4.000 214.520 295.600 215.920 ;
        RECT 4.000 213.880 296.000 214.520 ;
        RECT 4.000 212.480 295.600 213.880 ;
        RECT 4.000 211.160 296.000 212.480 ;
        RECT 4.000 209.760 295.600 211.160 ;
        RECT 4.000 209.120 296.000 209.760 ;
        RECT 4.000 207.720 295.600 209.120 ;
        RECT 4.000 206.400 296.000 207.720 ;
        RECT 4.000 205.000 295.600 206.400 ;
        RECT 4.000 204.360 296.000 205.000 ;
        RECT 4.000 202.960 295.600 204.360 ;
        RECT 4.000 202.320 296.000 202.960 ;
        RECT 4.000 200.920 295.600 202.320 ;
        RECT 4.000 199.600 296.000 200.920 ;
        RECT 4.000 198.200 295.600 199.600 ;
        RECT 4.000 197.560 296.000 198.200 ;
        RECT 4.000 196.160 295.600 197.560 ;
        RECT 4.000 194.840 296.000 196.160 ;
        RECT 4.000 193.440 295.600 194.840 ;
        RECT 4.000 192.800 296.000 193.440 ;
        RECT 4.000 191.400 295.600 192.800 ;
        RECT 4.000 190.760 296.000 191.400 ;
        RECT 4.000 189.360 295.600 190.760 ;
        RECT 4.000 188.040 296.000 189.360 ;
        RECT 4.000 186.640 295.600 188.040 ;
        RECT 4.000 186.000 296.000 186.640 ;
        RECT 4.000 184.600 295.600 186.000 ;
        RECT 4.000 183.280 296.000 184.600 ;
        RECT 4.000 181.880 295.600 183.280 ;
        RECT 4.000 181.240 296.000 181.880 ;
        RECT 4.000 179.840 295.600 181.240 ;
        RECT 4.000 179.200 296.000 179.840 ;
        RECT 4.000 177.800 295.600 179.200 ;
        RECT 4.000 176.480 296.000 177.800 ;
        RECT 4.000 175.080 295.600 176.480 ;
        RECT 4.000 174.440 296.000 175.080 ;
        RECT 4.000 173.040 295.600 174.440 ;
        RECT 4.000 172.400 296.000 173.040 ;
        RECT 4.000 171.000 295.600 172.400 ;
        RECT 4.000 169.680 296.000 171.000 ;
        RECT 4.000 168.280 295.600 169.680 ;
        RECT 4.000 167.640 296.000 168.280 ;
        RECT 4.000 166.240 295.600 167.640 ;
        RECT 4.000 164.920 296.000 166.240 ;
        RECT 4.000 163.520 295.600 164.920 ;
        RECT 4.000 162.880 296.000 163.520 ;
        RECT 4.000 161.480 295.600 162.880 ;
        RECT 4.000 160.840 296.000 161.480 ;
        RECT 4.000 159.440 295.600 160.840 ;
        RECT 4.000 158.120 296.000 159.440 ;
        RECT 4.000 156.720 295.600 158.120 ;
        RECT 4.000 156.080 296.000 156.720 ;
        RECT 4.000 154.680 295.600 156.080 ;
        RECT 4.000 153.360 296.000 154.680 ;
        RECT 4.000 151.960 295.600 153.360 ;
        RECT 4.000 151.320 296.000 151.960 ;
        RECT 4.000 149.920 295.600 151.320 ;
        RECT 4.000 149.280 296.000 149.920 ;
        RECT 4.000 147.880 295.600 149.280 ;
        RECT 4.000 146.560 296.000 147.880 ;
        RECT 4.000 145.160 295.600 146.560 ;
        RECT 4.000 144.520 296.000 145.160 ;
        RECT 4.000 143.120 295.600 144.520 ;
        RECT 4.000 141.800 296.000 143.120 ;
        RECT 4.000 140.400 295.600 141.800 ;
        RECT 4.000 139.760 296.000 140.400 ;
        RECT 4.000 138.360 295.600 139.760 ;
        RECT 4.000 137.720 296.000 138.360 ;
        RECT 4.000 136.320 295.600 137.720 ;
        RECT 4.000 135.000 296.000 136.320 ;
        RECT 4.000 133.600 295.600 135.000 ;
        RECT 4.000 132.960 296.000 133.600 ;
        RECT 4.000 131.560 295.600 132.960 ;
        RECT 4.000 130.240 296.000 131.560 ;
        RECT 4.000 128.840 295.600 130.240 ;
        RECT 4.000 128.200 296.000 128.840 ;
        RECT 4.000 126.800 295.600 128.200 ;
        RECT 4.000 126.160 296.000 126.800 ;
        RECT 4.000 124.760 295.600 126.160 ;
        RECT 4.000 123.440 296.000 124.760 ;
        RECT 4.000 122.040 295.600 123.440 ;
        RECT 4.000 121.400 296.000 122.040 ;
        RECT 4.000 120.000 295.600 121.400 ;
        RECT 4.000 119.360 296.000 120.000 ;
        RECT 4.000 117.960 295.600 119.360 ;
        RECT 4.000 116.640 296.000 117.960 ;
        RECT 4.000 115.240 295.600 116.640 ;
        RECT 4.000 114.600 296.000 115.240 ;
        RECT 4.000 113.200 295.600 114.600 ;
        RECT 4.000 111.880 296.000 113.200 ;
        RECT 4.000 110.480 295.600 111.880 ;
        RECT 4.000 109.840 296.000 110.480 ;
        RECT 4.000 108.440 295.600 109.840 ;
        RECT 4.000 107.800 296.000 108.440 ;
        RECT 4.000 106.400 295.600 107.800 ;
        RECT 4.000 105.080 296.000 106.400 ;
        RECT 4.000 103.680 295.600 105.080 ;
        RECT 4.000 103.040 296.000 103.680 ;
        RECT 4.000 101.640 295.600 103.040 ;
        RECT 4.000 100.320 296.000 101.640 ;
        RECT 4.000 98.920 295.600 100.320 ;
        RECT 4.000 98.280 296.000 98.920 ;
        RECT 4.000 96.880 295.600 98.280 ;
        RECT 4.000 96.240 296.000 96.880 ;
        RECT 4.000 94.840 295.600 96.240 ;
        RECT 4.000 93.520 296.000 94.840 ;
        RECT 4.000 92.120 295.600 93.520 ;
        RECT 4.000 91.480 296.000 92.120 ;
        RECT 4.000 90.080 295.600 91.480 ;
        RECT 4.000 88.760 296.000 90.080 ;
        RECT 4.000 87.360 295.600 88.760 ;
        RECT 4.000 86.720 296.000 87.360 ;
        RECT 4.000 85.320 295.600 86.720 ;
        RECT 4.000 84.680 296.000 85.320 ;
        RECT 4.000 83.280 295.600 84.680 ;
        RECT 4.000 81.960 296.000 83.280 ;
        RECT 4.000 80.560 295.600 81.960 ;
        RECT 4.000 79.920 296.000 80.560 ;
        RECT 4.000 78.520 295.600 79.920 ;
        RECT 4.000 77.200 296.000 78.520 ;
        RECT 4.000 75.840 295.600 77.200 ;
        RECT 4.400 75.800 295.600 75.840 ;
        RECT 4.400 75.160 296.000 75.800 ;
        RECT 4.400 74.440 295.600 75.160 ;
        RECT 4.000 73.760 295.600 74.440 ;
        RECT 4.000 73.120 296.000 73.760 ;
        RECT 4.000 71.720 295.600 73.120 ;
        RECT 4.000 70.400 296.000 71.720 ;
        RECT 4.000 69.000 295.600 70.400 ;
        RECT 4.000 68.360 296.000 69.000 ;
        RECT 4.000 66.960 295.600 68.360 ;
        RECT 4.000 65.640 296.000 66.960 ;
        RECT 4.000 64.240 295.600 65.640 ;
        RECT 4.000 63.600 296.000 64.240 ;
        RECT 4.000 62.200 295.600 63.600 ;
        RECT 4.000 61.560 296.000 62.200 ;
        RECT 4.000 60.160 295.600 61.560 ;
        RECT 4.000 58.840 296.000 60.160 ;
        RECT 4.000 57.440 295.600 58.840 ;
        RECT 4.000 56.800 296.000 57.440 ;
        RECT 4.000 55.400 295.600 56.800 ;
        RECT 4.000 54.760 296.000 55.400 ;
        RECT 4.000 53.360 295.600 54.760 ;
        RECT 4.000 52.040 296.000 53.360 ;
        RECT 4.000 50.640 295.600 52.040 ;
        RECT 4.000 50.000 296.000 50.640 ;
        RECT 4.000 48.600 295.600 50.000 ;
        RECT 4.000 47.280 296.000 48.600 ;
        RECT 4.000 45.880 295.600 47.280 ;
        RECT 4.000 45.240 296.000 45.880 ;
        RECT 4.000 43.840 295.600 45.240 ;
        RECT 4.000 43.200 296.000 43.840 ;
        RECT 4.000 41.800 295.600 43.200 ;
        RECT 4.000 40.480 296.000 41.800 ;
        RECT 4.000 39.080 295.600 40.480 ;
        RECT 4.000 38.440 296.000 39.080 ;
        RECT 4.000 37.040 295.600 38.440 ;
        RECT 4.000 35.720 296.000 37.040 ;
        RECT 4.000 34.320 295.600 35.720 ;
        RECT 4.000 33.680 296.000 34.320 ;
        RECT 4.000 32.280 295.600 33.680 ;
        RECT 4.000 31.640 296.000 32.280 ;
        RECT 4.000 30.240 295.600 31.640 ;
        RECT 4.000 28.920 296.000 30.240 ;
        RECT 4.000 27.520 295.600 28.920 ;
        RECT 4.000 26.880 296.000 27.520 ;
        RECT 4.000 25.480 295.600 26.880 ;
        RECT 4.000 24.160 296.000 25.480 ;
        RECT 4.000 22.760 295.600 24.160 ;
        RECT 4.000 22.120 296.000 22.760 ;
        RECT 4.000 20.720 295.600 22.120 ;
        RECT 4.000 20.080 296.000 20.720 ;
        RECT 4.000 18.680 295.600 20.080 ;
        RECT 4.000 17.360 296.000 18.680 ;
        RECT 4.000 15.960 295.600 17.360 ;
        RECT 4.000 15.320 296.000 15.960 ;
        RECT 4.000 13.920 295.600 15.320 ;
        RECT 4.000 12.600 296.000 13.920 ;
        RECT 4.000 11.200 295.600 12.600 ;
        RECT 4.000 10.560 296.000 11.200 ;
        RECT 4.000 9.160 295.600 10.560 ;
        RECT 4.000 8.520 296.000 9.160 ;
        RECT 4.000 7.120 295.600 8.520 ;
        RECT 4.000 5.800 296.000 7.120 ;
        RECT 4.000 4.400 295.600 5.800 ;
        RECT 4.000 3.760 296.000 4.400 ;
        RECT 4.000 2.360 295.600 3.760 ;
        RECT 4.000 1.720 296.000 2.360 ;
        RECT 4.000 0.855 295.600 1.720 ;
      LAYER met4 ;
        RECT 279.055 269.455 279.385 273.865 ;
  END
END spm_top
END LIBRARY

