

module __DESIGN__UNDER__TEST__
(
  mc,
  mp,
  clk,
  rst,
  prod,
  start,
  done,
  sin,
  shift,
  sout,
  tck,
  test
);

  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire \__BoundaryScanRegister_input_0__.dout ;
  wire \__BoundaryScanRegister_input_0__.sout ;
  wire \__BoundaryScanRegister_input_10__.dout ;
  wire \__BoundaryScanRegister_input_10__.sin ;
  wire \__BoundaryScanRegister_input_10__.sout ;
  wire \__BoundaryScanRegister_input_11__.dout ;
  wire \__BoundaryScanRegister_input_11__.sout ;
  wire \__BoundaryScanRegister_input_12__.dout ;
  wire \__BoundaryScanRegister_input_12__.sout ;
  wire \__BoundaryScanRegister_input_13__.dout ;
  wire \__BoundaryScanRegister_input_13__.sout ;
  wire \__BoundaryScanRegister_input_14__.dout ;
  wire \__BoundaryScanRegister_input_14__.sout ;
  wire \__BoundaryScanRegister_input_15__.dout ;
  wire \__BoundaryScanRegister_input_15__.sout ;
  wire \__BoundaryScanRegister_input_16__.dout ;
  wire \__BoundaryScanRegister_input_16__.sout ;
  wire \__BoundaryScanRegister_input_17__.dout ;
  wire \__BoundaryScanRegister_input_17__.sout ;
  wire \__BoundaryScanRegister_input_18__.dout ;
  wire \__BoundaryScanRegister_input_18__.sout ;
  wire \__BoundaryScanRegister_input_19__.dout ;
  wire \__BoundaryScanRegister_input_19__.sout ;
  wire \__BoundaryScanRegister_input_1__.dout ;
  wire \__BoundaryScanRegister_input_1__.sout ;
  wire \__BoundaryScanRegister_input_20__.dout ;
  wire \__BoundaryScanRegister_input_20__.sout ;
  wire \__BoundaryScanRegister_input_21__.dout ;
  wire \__BoundaryScanRegister_input_21__.sout ;
  wire \__BoundaryScanRegister_input_22__.dout ;
  wire \__BoundaryScanRegister_input_22__.sout ;
  wire \__BoundaryScanRegister_input_23__.dout ;
  wire \__BoundaryScanRegister_input_23__.sout ;
  wire \__BoundaryScanRegister_input_24__.dout ;
  wire \__BoundaryScanRegister_input_24__.sout ;
  wire \__BoundaryScanRegister_input_25__.dout ;
  wire \__BoundaryScanRegister_input_25__.sout ;
  wire \__BoundaryScanRegister_input_26__.dout ;
  wire \__BoundaryScanRegister_input_26__.sout ;
  wire \__BoundaryScanRegister_input_27__.dout ;
  wire \__BoundaryScanRegister_input_27__.sout ;
  wire \__BoundaryScanRegister_input_28__.dout ;
  wire \__BoundaryScanRegister_input_28__.sout ;
  wire \__BoundaryScanRegister_input_29__.dout ;
  wire \__BoundaryScanRegister_input_29__.sout ;
  wire \__BoundaryScanRegister_input_2__.dout ;
  wire \__BoundaryScanRegister_input_2__.sout ;
  wire \__BoundaryScanRegister_input_30__.dout ;
  wire \__BoundaryScanRegister_input_30__.sout ;
  wire \__BoundaryScanRegister_input_31__.dout ;
  wire \__BoundaryScanRegister_input_31__.sout ;
  wire \__BoundaryScanRegister_input_32__.dout ;
  wire \__BoundaryScanRegister_input_32__.sout ;
  wire \__BoundaryScanRegister_input_33__.dout ;
  wire \__BoundaryScanRegister_input_33__.sout ;
  wire \__BoundaryScanRegister_input_34__.dout ;
  wire \__BoundaryScanRegister_input_34__.sout ;
  wire \__BoundaryScanRegister_input_35__.dout ;
  wire \__BoundaryScanRegister_input_35__.sout ;
  wire \__BoundaryScanRegister_input_36__.dout ;
  wire \__BoundaryScanRegister_input_36__.sout ;
  wire \__BoundaryScanRegister_input_37__.dout ;
  wire \__BoundaryScanRegister_input_37__.sout ;
  wire \__BoundaryScanRegister_input_38__.dout ;
  wire \__BoundaryScanRegister_input_38__.sout ;
  wire \__BoundaryScanRegister_input_39__.dout ;
  wire \__BoundaryScanRegister_input_39__.sout ;
  wire \__BoundaryScanRegister_input_3__.dout ;
  wire \__BoundaryScanRegister_input_3__.sout ;
  wire \__BoundaryScanRegister_input_40__.dout ;
  wire \__BoundaryScanRegister_input_40__.sout ;
  wire \__BoundaryScanRegister_input_41__.dout ;
  wire \__BoundaryScanRegister_input_41__.sout ;
  wire \__BoundaryScanRegister_input_42__.dout ;
  wire \__BoundaryScanRegister_input_42__.sout ;
  wire \__BoundaryScanRegister_input_43__.dout ;
  wire \__BoundaryScanRegister_input_43__.sout ;
  wire \__BoundaryScanRegister_input_44__.dout ;
  wire \__BoundaryScanRegister_input_44__.sout ;
  wire \__BoundaryScanRegister_input_45__.dout ;
  wire \__BoundaryScanRegister_input_45__.sout ;
  wire \__BoundaryScanRegister_input_46__.dout ;
  wire \__BoundaryScanRegister_input_46__.sout ;
  wire \__BoundaryScanRegister_input_47__.dout ;
  wire \__BoundaryScanRegister_input_47__.sout ;
  wire \__BoundaryScanRegister_input_48__.dout ;
  wire \__BoundaryScanRegister_input_48__.sout ;
  wire \__BoundaryScanRegister_input_49__.dout ;
  wire \__BoundaryScanRegister_input_49__.sout ;
  wire \__BoundaryScanRegister_input_4__.dout ;
  wire \__BoundaryScanRegister_input_4__.sout ;
  wire \__BoundaryScanRegister_input_50__.dout ;
  wire \__BoundaryScanRegister_input_50__.sout ;
  wire \__BoundaryScanRegister_input_51__.dout ;
  wire \__BoundaryScanRegister_input_51__.sout ;
  wire \__BoundaryScanRegister_input_52__.dout ;
  wire \__BoundaryScanRegister_input_52__.sout ;
  wire \__BoundaryScanRegister_input_53__.dout ;
  wire \__BoundaryScanRegister_input_53__.sout ;
  wire \__BoundaryScanRegister_input_54__.dout ;
  wire \__BoundaryScanRegister_input_54__.sout ;
  wire \__BoundaryScanRegister_input_55__.dout ;
  wire \__BoundaryScanRegister_input_55__.sout ;
  wire \__BoundaryScanRegister_input_56__.dout ;
  wire \__BoundaryScanRegister_input_56__.sout ;
  wire \__BoundaryScanRegister_input_57__.dout ;
  wire \__BoundaryScanRegister_input_57__.sout ;
  wire \__BoundaryScanRegister_input_58__.dout ;
  wire \__BoundaryScanRegister_input_58__.sout ;
  wire \__BoundaryScanRegister_input_59__.dout ;
  wire \__BoundaryScanRegister_input_59__.sout ;
  wire \__BoundaryScanRegister_input_5__.dout ;
  wire \__BoundaryScanRegister_input_5__.sout ;
  wire \__BoundaryScanRegister_input_60__.dout ;
  wire \__BoundaryScanRegister_input_60__.sout ;
  wire \__BoundaryScanRegister_input_61__.dout ;
  wire \__BoundaryScanRegister_input_61__.sout ;
  wire \__BoundaryScanRegister_input_62__.dout ;
  wire \__BoundaryScanRegister_input_62__.sout ;
  wire \__BoundaryScanRegister_input_63__.dout ;
  wire \__BoundaryScanRegister_input_63__.sout ;
  wire \__BoundaryScanRegister_input_64__.dout ;
  wire \__BoundaryScanRegister_input_64__.sout ;
  wire \__BoundaryScanRegister_input_6__.dout ;
  wire \__BoundaryScanRegister_input_6__.sout ;
  wire \__BoundaryScanRegister_input_7__.dout ;
  wire \__BoundaryScanRegister_input_7__.sout ;
  wire \__BoundaryScanRegister_input_8__.dout ;
  wire \__BoundaryScanRegister_input_8__.sout ;
  wire \__BoundaryScanRegister_input_9__.dout ;
  wire \__BoundaryScanRegister_output_100__.sin ;
  wire \__BoundaryScanRegister_output_100__.sout ;
  wire \__BoundaryScanRegister_output_101__.sout ;
  wire \__BoundaryScanRegister_output_102__.sout ;
  wire \__BoundaryScanRegister_output_103__.sout ;
  wire \__BoundaryScanRegister_output_104__.sout ;
  wire \__BoundaryScanRegister_output_105__.sout ;
  wire \__BoundaryScanRegister_output_106__.sout ;
  wire \__BoundaryScanRegister_output_107__.sout ;
  wire \__BoundaryScanRegister_output_108__.sout ;
  wire \__BoundaryScanRegister_output_109__.sout ;
  wire \__BoundaryScanRegister_output_110__.sout ;
  wire \__BoundaryScanRegister_output_111__.sout ;
  wire \__BoundaryScanRegister_output_112__.sout ;
  wire \__BoundaryScanRegister_output_113__.sout ;
  wire \__BoundaryScanRegister_output_114__.sout ;
  wire \__BoundaryScanRegister_output_115__.sout ;
  wire \__BoundaryScanRegister_output_116__.sout ;
  wire \__BoundaryScanRegister_output_117__.sout ;
  wire \__BoundaryScanRegister_output_118__.sout ;
  wire \__BoundaryScanRegister_output_119__.sout ;
  wire \__BoundaryScanRegister_output_120__.sout ;
  wire \__BoundaryScanRegister_output_121__.sout ;
  wire \__BoundaryScanRegister_output_122__.sout ;
  wire \__BoundaryScanRegister_output_123__.sout ;
  wire \__BoundaryScanRegister_output_124__.sout ;
  wire \__BoundaryScanRegister_output_125__.sout ;
  wire \__BoundaryScanRegister_output_126__.sout ;
  wire \__BoundaryScanRegister_output_127__.sout ;
  wire \__BoundaryScanRegister_output_128__.sout ;
  wire \__BoundaryScanRegister_output_65__.sin ;
  wire \__BoundaryScanRegister_output_65__.sout ;
  wire \__BoundaryScanRegister_output_66__.sout ;
  wire \__BoundaryScanRegister_output_67__.sout ;
  wire \__BoundaryScanRegister_output_68__.sout ;
  wire \__BoundaryScanRegister_output_69__.sout ;
  wire \__BoundaryScanRegister_output_70__.sout ;
  wire \__BoundaryScanRegister_output_71__.sout ;
  wire \__BoundaryScanRegister_output_72__.sout ;
  wire \__BoundaryScanRegister_output_73__.sout ;
  wire \__BoundaryScanRegister_output_74__.sout ;
  wire \__BoundaryScanRegister_output_75__.sout ;
  wire \__BoundaryScanRegister_output_76__.sout ;
  wire \__BoundaryScanRegister_output_77__.sout ;
  wire \__BoundaryScanRegister_output_78__.sout ;
  wire \__BoundaryScanRegister_output_79__.sout ;
  wire \__BoundaryScanRegister_output_80__.sout ;
  wire \__BoundaryScanRegister_output_81__.sout ;
  wire \__BoundaryScanRegister_output_82__.sout ;
  wire \__BoundaryScanRegister_output_83__.sout ;
  wire \__BoundaryScanRegister_output_84__.sout ;
  wire \__BoundaryScanRegister_output_85__.sout ;
  wire \__BoundaryScanRegister_output_86__.sout ;
  wire \__BoundaryScanRegister_output_87__.sout ;
  wire \__BoundaryScanRegister_output_88__.sout ;
  wire \__BoundaryScanRegister_output_89__.sout ;
  wire \__BoundaryScanRegister_output_90__.sout ;
  wire \__BoundaryScanRegister_output_91__.sout ;
  wire \__BoundaryScanRegister_output_92__.sout ;
  wire \__BoundaryScanRegister_output_93__.sout ;
  wire \__BoundaryScanRegister_output_94__.sout ;
  wire \__BoundaryScanRegister_output_95__.sout ;
  wire \__BoundaryScanRegister_output_96__.sout ;
  wire \__BoundaryScanRegister_output_97__.sout ;
  wire \__BoundaryScanRegister_output_98__.sout ;
  wire \__uuf__._0000_ ;
  wire \__uuf__._0001_ ;
  wire \__uuf__._0002_ ;
  wire \__uuf__._0003_ ;
  wire \__uuf__._0004_ ;
  wire \__uuf__._0005_ ;
  wire \__uuf__._0006_ ;
  wire \__uuf__._0007_ ;
  wire \__uuf__._0008_ ;
  wire \__uuf__._0009_ ;
  wire \__uuf__._0010_ ;
  wire \__uuf__._0011_ ;
  wire \__uuf__._0012_ ;
  wire \__uuf__._0013_ ;
  wire \__uuf__._0014_ ;
  wire \__uuf__._0015_ ;
  wire \__uuf__._0016_ ;
  wire \__uuf__._0017_ ;
  wire \__uuf__._0018_ ;
  wire \__uuf__._0019_ ;
  wire \__uuf__._0020_ ;
  wire \__uuf__._0021_ ;
  wire \__uuf__._0022_ ;
  wire \__uuf__._0023_ ;
  wire \__uuf__._0024_ ;
  wire \__uuf__._0025_ ;
  wire \__uuf__._0026_ ;
  wire \__uuf__._0027_ ;
  wire \__uuf__._0028_ ;
  wire \__uuf__._0029_ ;
  wire \__uuf__._0030_ ;
  wire \__uuf__._0031_ ;
  wire \__uuf__._0032_ ;
  wire \__uuf__._0033_ ;
  wire \__uuf__._0034_ ;
  wire \__uuf__._0035_ ;
  wire \__uuf__._0036_ ;
  wire \__uuf__._0037_ ;
  wire \__uuf__._0038_ ;
  wire \__uuf__._0039_ ;
  wire \__uuf__._0040_ ;
  wire \__uuf__._0041_ ;
  wire \__uuf__._0042_ ;
  wire \__uuf__._0043_ ;
  wire \__uuf__._0044_ ;
  wire \__uuf__._0045_ ;
  wire \__uuf__._0046_ ;
  wire \__uuf__._0047_ ;
  wire \__uuf__._0048_ ;
  wire \__uuf__._0049_ ;
  wire \__uuf__._0050_ ;
  wire \__uuf__._0051_ ;
  wire \__uuf__._0052_ ;
  wire \__uuf__._0053_ ;
  wire \__uuf__._0054_ ;
  wire \__uuf__._0055_ ;
  wire \__uuf__._0056_ ;
  wire \__uuf__._0057_ ;
  wire \__uuf__._0058_ ;
  wire \__uuf__._0059_ ;
  wire \__uuf__._0060_ ;
  wire \__uuf__._0061_ ;
  wire \__uuf__._0062_ ;
  wire \__uuf__._0063_ ;
  wire \__uuf__._0064_ ;
  wire \__uuf__._0065_ ;
  wire \__uuf__._0066_ ;
  wire \__uuf__._0067_ ;
  wire \__uuf__._0068_ ;
  wire \__uuf__._0069_ ;
  wire \__uuf__._0070_ ;
  wire \__uuf__._0071_ ;
  wire \__uuf__._0072_ ;
  wire \__uuf__._0073_ ;
  wire \__uuf__._0074_ ;
  wire \__uuf__._0075_ ;
  wire \__uuf__._0076_ ;
  wire \__uuf__._0077_ ;
  wire \__uuf__._0078_ ;
  wire \__uuf__._0079_ ;
  wire \__uuf__._0080_ ;
  wire \__uuf__._0081_ ;
  wire \__uuf__._0082_ ;
  wire \__uuf__._0083_ ;
  wire \__uuf__._0084_ ;
  wire \__uuf__._0085_ ;
  wire \__uuf__._0086_ ;
  wire \__uuf__._0087_ ;
  wire \__uuf__._0088_ ;
  wire \__uuf__._0089_ ;
  wire \__uuf__._0090_ ;
  wire \__uuf__._0091_ ;
  wire \__uuf__._0092_ ;
  wire \__uuf__._0093_ ;
  wire \__uuf__._0094_ ;
  wire \__uuf__._0095_ ;
  wire \__uuf__._0096_ ;
  wire \__uuf__._0097_ ;
  wire \__uuf__._0098_ ;
  wire \__uuf__._0099_ ;
  wire \__uuf__._0100_ ;
  wire \__uuf__._0101_ ;
  wire \__uuf__._0102_ ;
  wire \__uuf__._0103_ ;
  wire \__uuf__._0104_ ;
  wire \__uuf__._0105_ ;
  wire \__uuf__._0106_ ;
  wire \__uuf__._0107_ ;
  wire \__uuf__._0108_ ;
  wire \__uuf__._0109_ ;
  wire \__uuf__._0110_ ;
  wire \__uuf__._0111_ ;
  wire \__uuf__._0112_ ;
  wire \__uuf__._0113_ ;
  wire \__uuf__._0114_ ;
  wire \__uuf__._0115_ ;
  wire \__uuf__._0116_ ;
  wire \__uuf__._0117_ ;
  wire \__uuf__._0118_ ;
  wire \__uuf__._0119_ ;
  wire \__uuf__._0120_ ;
  wire \__uuf__._0121_ ;
  wire \__uuf__._0122_ ;
  wire \__uuf__._0123_ ;
  wire \__uuf__._0124_ ;
  wire \__uuf__._0125_ ;
  wire \__uuf__._0126_ ;
  wire \__uuf__._0127_ ;
  wire \__uuf__._0128_ ;
  wire \__uuf__._0129_ ;
  wire \__uuf__._0130_ ;
  wire \__uuf__._0131_ ;
  wire \__uuf__._0132_ ;
  wire \__uuf__._0133_ ;
  wire \__uuf__._0134_ ;
  wire \__uuf__._0135_ ;
  wire \__uuf__._0136_ ;
  wire \__uuf__._0137_ ;
  wire \__uuf__._0138_ ;
  wire \__uuf__._0139_ ;
  wire \__uuf__._0140_ ;
  wire \__uuf__._0141_ ;
  wire \__uuf__._0142_ ;
  wire \__uuf__._0143_ ;
  wire \__uuf__._0144_ ;
  wire \__uuf__._0145_ ;
  wire \__uuf__._0146_ ;
  wire \__uuf__._0147_ ;
  wire \__uuf__._0148_ ;
  wire \__uuf__._0149_ ;
  wire \__uuf__._0150_ ;
  wire \__uuf__._0151_ ;
  wire \__uuf__._0152_ ;
  wire \__uuf__._0153_ ;
  wire \__uuf__._0154_ ;
  wire \__uuf__._0155_ ;
  wire \__uuf__._0156_ ;
  wire \__uuf__._0157_ ;
  wire \__uuf__._0158_ ;
  wire \__uuf__._0159_ ;
  wire \__uuf__._0160_ ;
  wire \__uuf__._0161_ ;
  wire \__uuf__._0162_ ;
  wire \__uuf__._0163_ ;
  wire \__uuf__._0164_ ;
  wire \__uuf__._0165_ ;
  wire \__uuf__._0166_ ;
  wire \__uuf__._0167_ ;
  wire \__uuf__._0168_ ;
  wire \__uuf__._0169_ ;
  wire \__uuf__._0170_ ;
  wire \__uuf__._0171_ ;
  wire \__uuf__._0172_ ;
  wire \__uuf__._0173_ ;
  wire \__uuf__._0174_ ;
  wire \__uuf__._0175_ ;
  wire \__uuf__._0176_ ;
  wire \__uuf__._0177_ ;
  wire \__uuf__._0178_ ;
  wire \__uuf__._0179_ ;
  wire \__uuf__._0180_ ;
  wire \__uuf__._0181_ ;
  wire \__uuf__._0182_ ;
  wire \__uuf__._0183_ ;
  wire \__uuf__._0184_ ;
  wire \__uuf__._0185_ ;
  wire \__uuf__._0186_ ;
  wire \__uuf__._0187_ ;
  wire \__uuf__._0188_ ;
  wire \__uuf__._0189_ ;
  wire \__uuf__._0190_ ;
  wire \__uuf__._0191_ ;
  wire \__uuf__._0192_ ;
  wire \__uuf__._0193_ ;
  wire \__uuf__._0194_ ;
  wire \__uuf__._0195_ ;
  wire \__uuf__._0196_ ;
  wire \__uuf__._0197_ ;
  wire \__uuf__._0198_ ;
  wire \__uuf__._0199_ ;
  wire \__uuf__._0200_ ;
  wire \__uuf__._0201_ ;
  wire \__uuf__._0202_ ;
  wire \__uuf__._0203_ ;
  wire \__uuf__._0204_ ;
  wire \__uuf__._0205_ ;
  wire \__uuf__._0206_ ;
  wire \__uuf__._0207_ ;
  wire \__uuf__._0208_ ;
  wire \__uuf__._0209_ ;
  wire \__uuf__._0210_ ;
  wire \__uuf__._0211_ ;
  wire \__uuf__._0212_ ;
  wire \__uuf__._0213_ ;
  wire \__uuf__._0214_ ;
  wire \__uuf__._0215_ ;
  wire \__uuf__._0216_ ;
  wire \__uuf__._0217_ ;
  wire \__uuf__._0218_ ;
  wire \__uuf__._0219_ ;
  wire \__uuf__._0220_ ;
  wire \__uuf__._0221_ ;
  wire \__uuf__._0222_ ;
  wire \__uuf__._0223_ ;
  wire \__uuf__._0224_ ;
  wire \__uuf__._0225_ ;
  wire \__uuf__._0226_ ;
  wire \__uuf__._0227_ ;
  wire \__uuf__._0228_ ;
  wire \__uuf__._0229_ ;
  wire \__uuf__._0230_ ;
  wire \__uuf__._0231_ ;
  wire \__uuf__._0232_ ;
  wire \__uuf__._0233_ ;
  wire \__uuf__._0234_ ;
  wire \__uuf__._0235_ ;
  wire \__uuf__._0236_ ;
  wire \__uuf__._0237_ ;
  wire \__uuf__._0238_ ;
  wire \__uuf__._0239_ ;
  wire \__uuf__._0240_ ;
  wire \__uuf__._0241_ ;
  wire \__uuf__._0242_ ;
  wire \__uuf__._0243_ ;
  wire \__uuf__._0244_ ;
  wire \__uuf__._0245_ ;
  wire \__uuf__._0246_ ;
  wire \__uuf__._0247_ ;
  wire \__uuf__._0248_ ;
  wire \__uuf__._0249_ ;
  wire \__uuf__._0250_ ;
  wire \__uuf__._0251_ ;
  wire \__uuf__._0252_ ;
  wire \__uuf__._0253_ ;
  wire \__uuf__._0254_ ;
  wire \__uuf__._0255_ ;
  wire \__uuf__._0256_ ;
  wire \__uuf__._0257_ ;
  wire \__uuf__._0258_ ;
  wire \__uuf__._0259_ ;
  wire \__uuf__._0260_ ;
  wire \__uuf__._0261_ ;
  wire \__uuf__._0262_ ;
  wire \__uuf__._0263_ ;
  wire \__uuf__._0264_ ;
  wire \__uuf__._0265_ ;
  wire \__uuf__._0266_ ;
  wire \__uuf__._0267_ ;
  wire \__uuf__._0268_ ;
  wire \__uuf__._0269_ ;
  wire \__uuf__._0270_ ;
  wire \__uuf__._0271_ ;
  wire \__uuf__._0272_ ;
  wire \__uuf__._0273_ ;
  wire \__uuf__._0274_ ;
  wire \__uuf__._0275_ ;
  wire \__uuf__._0276_ ;
  wire \__uuf__._0277_ ;
  wire \__uuf__._0278_ ;
  wire \__uuf__._0279_ ;
  wire \__uuf__._0280_ ;
  wire \__uuf__._0281_ ;
  wire \__uuf__._0282_ ;
  wire \__uuf__._0283_ ;
  wire \__uuf__._0284_ ;
  wire \__uuf__._0285_ ;
  wire \__uuf__._0286_ ;
  wire \__uuf__._0287_ ;
  wire \__uuf__._0288_ ;
  wire \__uuf__._0289_ ;
  wire \__uuf__._0290_ ;
  wire \__uuf__._0291_ ;
  wire \__uuf__._0292_ ;
  wire \__uuf__._0293_ ;
  wire \__uuf__._0294_ ;
  wire \__uuf__._0295_ ;
  wire \__uuf__._0296_ ;
  wire \__uuf__._0297_ ;
  wire \__uuf__._0298_ ;
  wire \__uuf__._0299_ ;
  wire \__uuf__._0300_ ;
  wire \__uuf__._0301_ ;
  wire \__uuf__._0302_ ;
  wire \__uuf__._0303_ ;
  wire \__uuf__._0304_ ;
  wire \__uuf__._0305_ ;
  wire \__uuf__._0306_ ;
  wire \__uuf__._0307_ ;
  wire \__uuf__._0308_ ;
  wire \__uuf__._0309_ ;
  wire \__uuf__._0310_ ;
  wire \__uuf__._0311_ ;
  wire \__uuf__._0312_ ;
  wire \__uuf__._0313_ ;
  wire \__uuf__._0314_ ;
  wire \__uuf__._0315_ ;
  wire \__uuf__._0316_ ;
  wire \__uuf__._0317_ ;
  wire \__uuf__._0318_ ;
  wire \__uuf__._0319_ ;
  wire \__uuf__._0320_ ;
  wire \__uuf__._0321_ ;
  wire \__uuf__._0322_ ;
  wire \__uuf__._0323_ ;
  wire \__uuf__._0324_ ;
  wire \__uuf__._0325_ ;
  wire \__uuf__._0326_ ;
  wire \__uuf__._0327_ ;
  wire \__uuf__._0328_ ;
  wire \__uuf__._0329_ ;
  wire \__uuf__._0330_ ;
  wire \__uuf__._0331_ ;
  wire \__uuf__._0332_ ;
  wire \__uuf__._0333_ ;
  wire \__uuf__._0334_ ;
  wire \__uuf__._0335_ ;
  wire \__uuf__._0336_ ;
  wire \__uuf__._0337_ ;
  wire \__uuf__._0338_ ;
  wire \__uuf__._0339_ ;
  wire \__uuf__._0340_ ;
  wire \__uuf__._0341_ ;
  wire \__uuf__._0342_ ;
  wire \__uuf__._0343_ ;
  wire \__uuf__._0344_ ;
  wire \__uuf__._0345_ ;
  wire \__uuf__._0346_ ;
  wire \__uuf__._0347_ ;
  wire \__uuf__._0348_ ;
  wire \__uuf__._0349_ ;
  wire \__uuf__._0350_ ;
  wire \__uuf__._0351_ ;
  wire \__uuf__._0352_ ;
  wire \__uuf__._0353_ ;
  wire \__uuf__._0354_ ;
  wire \__uuf__._0355_ ;
  wire \__uuf__._0356_ ;
  wire \__uuf__._0357_ ;
  wire \__uuf__._0358_ ;
  wire \__uuf__._0359_ ;
  wire \__uuf__._0360_ ;
  wire \__uuf__._0361_ ;
  wire \__uuf__._0362_ ;
  wire \__uuf__._0363_ ;
  wire \__uuf__._0364_ ;
  wire \__uuf__._0365_ ;
  wire \__uuf__._0366_ ;
  wire \__uuf__._0367_ ;
  wire \__uuf__._0368_ ;
  wire \__uuf__._0369_ ;
  wire \__uuf__._0370_ ;
  wire \__uuf__._0371_ ;
  wire \__uuf__._0372_ ;
  wire \__uuf__._0373_ ;
  wire \__uuf__._0374_ ;
  wire \__uuf__._0375_ ;
  wire \__uuf__._0376_ ;
  wire \__uuf__._0377_ ;
  wire \__uuf__._0378_ ;
  wire \__uuf__._0379_ ;
  wire \__uuf__._0380_ ;
  wire \__uuf__._0381_ ;
  wire \__uuf__._0382_ ;
  wire \__uuf__._0383_ ;
  wire \__uuf__._0384_ ;
  wire \__uuf__._0385_ ;
  wire \__uuf__._0386_ ;
  wire \__uuf__._0387_ ;
  wire \__uuf__._0388_ ;
  wire \__uuf__._0389_ ;
  wire \__uuf__._0390_ ;
  wire \__uuf__._0391_ ;
  wire \__uuf__._0392_ ;
  wire \__uuf__._0393_ ;
  wire \__uuf__._0394_ ;
  wire \__uuf__._0395_ ;
  wire \__uuf__._0396_ ;
  wire \__uuf__._0397_ ;
  wire \__uuf__._0398_ ;
  wire \__uuf__._0399_ ;
  wire \__uuf__._0400_ ;
  wire \__uuf__._0401_ ;
  wire \__uuf__._0402_ ;
  wire \__uuf__._0403_ ;
  wire \__uuf__._0404_ ;
  wire \__uuf__._0405_ ;
  wire \__uuf__._0406_ ;
  wire \__uuf__._0407_ ;
  wire \__uuf__._0408_ ;
  wire \__uuf__._0409_ ;
  wire \__uuf__._0410_ ;
  wire \__uuf__._0411_ ;
  wire \__uuf__._0412_ ;
  wire \__uuf__._0413_ ;
  wire \__uuf__._0414_ ;
  wire \__uuf__._0415_ ;
  wire \__uuf__._0416_ ;
  wire \__uuf__._0417_ ;
  wire \__uuf__._0418_ ;
  wire \__uuf__._0419_ ;
  wire \__uuf__._0420_ ;
  wire \__uuf__._0421_ ;
  wire \__uuf__._0422_ ;
  wire \__uuf__._0423_ ;
  wire \__uuf__._0424_ ;
  wire \__uuf__._0425_ ;
  wire \__uuf__._0426_ ;
  wire \__uuf__._0427_ ;
  wire \__uuf__._0428_ ;
  wire \__uuf__._0429_ ;
  wire \__uuf__._0430_ ;
  wire \__uuf__._0431_ ;
  wire \__uuf__._0432_ ;
  wire \__uuf__._0433_ ;
  wire \__uuf__._0434_ ;
  wire \__uuf__._0435_ ;
  wire \__uuf__._0436_ ;
  wire \__uuf__._0437_ ;
  wire \__uuf__._0438_ ;
  wire \__uuf__._0439_ ;
  wire \__uuf__._0440_ ;
  wire \__uuf__._0441_ ;
  wire \__uuf__._0442_ ;
  wire \__uuf__._0443_ ;
  wire \__uuf__._0444_ ;
  wire \__uuf__._0445_ ;
  wire \__uuf__._0446_ ;
  wire \__uuf__._0447_ ;
  wire \__uuf__._0448_ ;
  wire \__uuf__._0449_ ;
  wire \__uuf__._0450_ ;
  wire \__uuf__._0451_ ;
  wire \__uuf__._0452_ ;
  wire \__uuf__._0453_ ;
  wire \__uuf__._0454_ ;
  wire \__uuf__._0455_ ;
  wire \__uuf__._0456_ ;
  wire \__uuf__._0457_ ;
  wire \__uuf__._0458_ ;
  wire \__uuf__._0459_ ;
  wire \__uuf__._0460_ ;
  wire \__uuf__._0461_ ;
  wire \__uuf__._0462_ ;
  wire \__uuf__._0463_ ;
  wire \__uuf__._0464_ ;
  wire \__uuf__._0465_ ;
  wire \__uuf__._0466_ ;
  wire \__uuf__._0467_ ;
  wire \__uuf__._0468_ ;
  wire \__uuf__._0469_ ;
  wire \__uuf__._0470_ ;
  wire \__uuf__._0471_ ;
  wire \__uuf__._0472_ ;
  wire \__uuf__._0473_ ;
  wire \__uuf__._0474_ ;
  wire \__uuf__._0475_ ;
  wire \__uuf__._0476_ ;
  wire \__uuf__._0477_ ;
  wire \__uuf__._0478_ ;
  wire \__uuf__._0479_ ;
  wire \__uuf__._0480_ ;
  wire \__uuf__._0481_ ;
  wire \__uuf__._0482_ ;
  wire \__uuf__._0483_ ;
  wire \__uuf__._0484_ ;
  wire \__uuf__._0485_ ;
  wire \__uuf__._0486_ ;
  wire \__uuf__._0487_ ;
  wire \__uuf__._0488_ ;
  wire \__uuf__._0489_ ;
  wire \__uuf__._0490_ ;
  wire \__uuf__._0491_ ;
  wire \__uuf__._0492_ ;
  wire \__uuf__._0493_ ;
  wire \__uuf__._0494_ ;
  wire \__uuf__._0495_ ;
  wire \__uuf__._0496_ ;
  wire \__uuf__._0497_ ;
  wire \__uuf__._0498_ ;
  wire \__uuf__._0499_ ;
  wire \__uuf__._0500_ ;
  wire \__uuf__._0501_ ;
  wire \__uuf__._0502_ ;
  wire \__uuf__._0503_ ;
  wire \__uuf__._0504_ ;
  wire \__uuf__._0505_ ;
  wire \__uuf__._0506_ ;
  wire \__uuf__._0507_ ;
  wire \__uuf__._0508_ ;
  wire \__uuf__._0509_ ;
  wire \__uuf__._0510_ ;
  wire \__uuf__._0511_ ;
  wire \__uuf__._0512_ ;
  wire \__uuf__._0513_ ;
  wire \__uuf__._0514_ ;
  wire \__uuf__._0515_ ;
  wire \__uuf__._0516_ ;
  wire \__uuf__._0517_ ;
  wire \__uuf__._0518_ ;
  wire \__uuf__._0519_ ;
  wire \__uuf__._0520_ ;
  wire \__uuf__._0521_ ;
  wire \__uuf__._0522_ ;
  wire \__uuf__._0523_ ;
  wire \__uuf__._0524_ ;
  wire \__uuf__._0525_ ;
  wire \__uuf__._0526_ ;
  wire \__uuf__._0527_ ;
  wire \__uuf__._0528_ ;
  wire \__uuf__._0529_ ;
  wire \__uuf__._0530_ ;
  wire \__uuf__._0531_ ;
  wire \__uuf__._0532_ ;
  wire \__uuf__._0533_ ;
  wire \__uuf__._0534_ ;
  wire \__uuf__._0535_ ;
  wire \__uuf__._0536_ ;
  wire \__uuf__._0537_ ;
  wire \__uuf__._0538_ ;
  wire \__uuf__._0539_ ;
  wire \__uuf__._0540_ ;
  wire \__uuf__._0541_ ;
  wire \__uuf__._0542_ ;
  wire \__uuf__._0543_ ;
  wire \__uuf__._0544_ ;
  wire \__uuf__._0545_ ;
  wire \__uuf__._0546_ ;
  wire \__uuf__._0547_ ;
  wire \__uuf__._0548_ ;
  wire \__uuf__._0549_ ;
  wire \__uuf__._0550_ ;
  wire \__uuf__._0551_ ;
  wire \__uuf__._0552_ ;
  wire \__uuf__._0553_ ;
  wire \__uuf__._0554_ ;
  wire \__uuf__._0555_ ;
  wire \__uuf__._0556_ ;
  wire \__uuf__._0557_ ;
  wire \__uuf__._0558_ ;
  wire \__uuf__._0559_ ;
  wire \__uuf__._0560_ ;
  wire \__uuf__._0561_ ;
  wire \__uuf__._0562_ ;
  wire \__uuf__._0563_ ;
  wire \__uuf__._0564_ ;
  wire \__uuf__._0565_ ;
  wire \__uuf__._0566_ ;
  wire \__uuf__._0567_ ;
  wire \__uuf__._0568_ ;
  wire \__uuf__._0569_ ;
  wire \__uuf__._0570_ ;
  wire \__uuf__._0571_ ;
  wire \__uuf__._0572_ ;
  wire \__uuf__._0573_ ;
  wire \__uuf__._0574_ ;
  wire \__uuf__._0575_ ;
  wire \__uuf__._0576_ ;
  wire \__uuf__._0577_ ;
  wire \__uuf__._0578_ ;
  wire \__uuf__._0579_ ;
  wire \__uuf__._0580_ ;
  wire \__uuf__._0581_ ;
  wire \__uuf__._0582_ ;
  wire \__uuf__._0583_ ;
  wire \__uuf__._0584_ ;
  wire \__uuf__._0585_ ;
  wire \__uuf__._0586_ ;
  wire \__uuf__._0587_ ;
  wire \__uuf__._0588_ ;
  wire \__uuf__._0589_ ;
  wire \__uuf__._0590_ ;
  wire \__uuf__._0591_ ;
  wire \__uuf__._0592_ ;
  wire \__uuf__._0593_ ;
  wire \__uuf__._0594_ ;
  wire \__uuf__._0595_ ;
  wire \__uuf__._0596_ ;
  wire \__uuf__._0597_ ;
  wire \__uuf__._0598_ ;
  wire \__uuf__._0599_ ;
  wire \__uuf__._0600_ ;
  wire \__uuf__._0601_ ;
  wire \__uuf__._0602_ ;
  wire \__uuf__._0603_ ;
  wire \__uuf__._0604_ ;
  wire \__uuf__._0605_ ;
  wire \__uuf__._0606_ ;
  wire \__uuf__._0607_ ;
  wire \__uuf__._0608_ ;
  wire \__uuf__._0609_ ;
  wire \__uuf__._0610_ ;
  wire \__uuf__._0611_ ;
  wire \__uuf__._0612_ ;
  wire \__uuf__._0613_ ;
  wire \__uuf__._0614_ ;
  wire \__uuf__._0615_ ;
  wire \__uuf__._0616_ ;
  wire \__uuf__._0617_ ;
  wire \__uuf__._0618_ ;
  wire \__uuf__._0619_ ;
  wire \__uuf__._0620_ ;
  wire \__uuf__._0621_ ;
  wire \__uuf__._0622_ ;
  wire \__uuf__._0623_ ;
  wire \__uuf__._0624_ ;
  wire \__uuf__._0625_ ;
  wire \__uuf__._0626_ ;
  wire \__uuf__._0627_ ;
  wire \__uuf__._0628_ ;
  wire \__uuf__._0629_ ;
  wire \__uuf__._0630_ ;
  wire \__uuf__._0631_ ;
  wire \__uuf__._0632_ ;
  wire \__uuf__._0633_ ;
  wire \__uuf__._0634_ ;
  wire \__uuf__._0635_ ;
  wire \__uuf__._0636_ ;
  wire \__uuf__._0637_ ;
  wire \__uuf__._0638_ ;
  wire \__uuf__._0639_ ;
  wire \__uuf__._0640_ ;
  wire \__uuf__._0641_ ;
  wire \__uuf__._0642_ ;
  wire \__uuf__._0643_ ;
  wire \__uuf__._0644_ ;
  wire \__uuf__._0645_ ;
  wire \__uuf__._0646_ ;
  wire \__uuf__._0647_ ;
  wire \__uuf__._0648_ ;
  wire \__uuf__._0649_ ;
  wire \__uuf__._0650_ ;
  wire \__uuf__._0651_ ;
  wire \__uuf__._0652_ ;
  wire \__uuf__._0653_ ;
  wire \__uuf__._0654_ ;
  wire \__uuf__._0655_ ;
  wire \__uuf__._0656_ ;
  wire \__uuf__._0657_ ;
  wire \__uuf__._0658_ ;
  wire \__uuf__._0659_ ;
  wire \__uuf__._0660_ ;
  wire \__uuf__._0661_ ;
  wire \__uuf__._0662_ ;
  wire \__uuf__._0663_ ;
  wire \__uuf__._0664_ ;
  wire \__uuf__._0665_ ;
  wire \__uuf__._0666_ ;
  wire \__uuf__._0667_ ;
  wire \__uuf__._0668_ ;
  wire \__uuf__._0669_ ;
  wire \__uuf__._0670_ ;
  wire \__uuf__._0671_ ;
  wire \__uuf__._0672_ ;
  wire \__uuf__._0673_ ;
  wire \__uuf__._0674_ ;
  wire \__uuf__._0675_ ;
  wire \__uuf__._0676_ ;
  wire \__uuf__._0677_ ;
  wire \__uuf__._0678_ ;
  wire \__uuf__._0679_ ;
  wire \__uuf__._0680_ ;
  wire \__uuf__._0681_ ;
  wire \__uuf__._0682_ ;
  wire \__uuf__._0683_ ;
  wire \__uuf__._0684_ ;
  wire \__uuf__._0685_ ;
  wire \__uuf__._0686_ ;
  wire \__uuf__._0687_ ;
  wire \__uuf__._0688_ ;
  wire \__uuf__._0689_ ;
  wire \__uuf__._0690_ ;
  wire \__uuf__._0691_ ;
  wire \__uuf__._0692_ ;
  wire \__uuf__._0693_ ;
  wire \__uuf__._0694_ ;
  wire \__uuf__._0695_ ;
  wire \__uuf__._0696_ ;
  wire \__uuf__._0697_ ;
  wire \__uuf__._0698_ ;
  wire \__uuf__._0699_ ;
  wire \__uuf__._0700_ ;
  wire \__uuf__._0701_ ;
  wire \__uuf__._0702_ ;
  wire \__uuf__._0703_ ;
  wire \__uuf__._0704_ ;
  wire \__uuf__._0705_ ;
  wire \__uuf__._0706_ ;
  wire \__uuf__._0707_ ;
  wire \__uuf__._0708_ ;
  wire \__uuf__._0709_ ;
  wire \__uuf__._0710_ ;
  wire \__uuf__._0711_ ;
  wire \__uuf__._0712_ ;
  wire \__uuf__._0713_ ;
  wire \__uuf__._0714_ ;
  wire \__uuf__._0715_ ;
  wire \__uuf__._0716_ ;
  wire \__uuf__._0717_ ;
  wire \__uuf__._0718_ ;
  wire \__uuf__._0719_ ;
  wire \__uuf__._0720_ ;
  wire \__uuf__._0721_ ;
  wire \__uuf__._0722_ ;
  wire \__uuf__._0723_ ;
  wire \__uuf__._0724_ ;
  wire \__uuf__._0725_ ;
  wire \__uuf__._0726_ ;
  wire \__uuf__._0727_ ;
  wire \__uuf__._0728_ ;
  wire \__uuf__._0729_ ;
  wire \__uuf__._0730_ ;
  wire \__uuf__._0731_ ;
  wire \__uuf__._0732_ ;
  wire \__uuf__._0733_ ;
  wire \__uuf__._0734_ ;
  wire \__uuf__._0735_ ;
  wire \__uuf__._0736_ ;
  wire \__uuf__._0737_ ;
  wire \__uuf__._0738_ ;
  wire \__uuf__._0739_ ;
  wire \__uuf__._0740_ ;
  wire \__uuf__._0741_ ;
  wire \__uuf__._0742_ ;
  wire \__uuf__._0743_ ;
  wire \__uuf__._0744_ ;
  wire \__uuf__._0745_ ;
  wire \__uuf__._0746_ ;
  wire \__uuf__._0747_ ;
  wire \__uuf__._0748_ ;
  wire \__uuf__._0749_ ;
  wire \__uuf__._0750_ ;
  wire \__uuf__._0751_ ;
  wire \__uuf__._0752_ ;
  wire \__uuf__._0753_ ;
  wire \__uuf__._0754_ ;
  wire \__uuf__._0755_ ;
  wire \__uuf__._0756_ ;
  wire \__uuf__._0757_ ;
  wire \__uuf__._0758_ ;
  wire \__uuf__._0759_ ;
  wire \__uuf__._0760_ ;
  wire \__uuf__._0761_ ;
  wire \__uuf__._0762_ ;
  wire \__uuf__._0763_ ;
  wire \__uuf__._0764_ ;
  wire \__uuf__._0765_ ;
  wire \__uuf__._0766_ ;
  wire \__uuf__._0767_ ;
  wire \__uuf__._0768_ ;
  wire \__uuf__._0769_ ;
  wire \__uuf__._0770_ ;
  wire \__uuf__._0771_ ;
  wire \__uuf__._0772_ ;
  wire \__uuf__._0773_ ;
  wire \__uuf__._0774_ ;
  wire \__uuf__._0775_ ;
  wire \__uuf__._0776_ ;
  wire \__uuf__._0777_ ;
  wire \__uuf__._0778_ ;
  wire \__uuf__._0779_ ;
  wire \__uuf__._0780_ ;
  wire \__uuf__._0781_ ;
  wire \__uuf__._0782_ ;
  wire \__uuf__._0783_ ;
  wire \__uuf__._0784_ ;
  wire \__uuf__._0785_ ;
  wire \__uuf__._0786_ ;
  wire \__uuf__._0787_ ;
  wire \__uuf__._0788_ ;
  wire \__uuf__._0789_ ;
  wire \__uuf__._0790_ ;
  wire \__uuf__._0791_ ;
  wire \__uuf__._0792_ ;
  wire \__uuf__._0793_ ;
  wire \__uuf__._0794_ ;
  wire \__uuf__._0795_ ;
  wire \__uuf__._0796_ ;
  wire \__uuf__._0797_ ;
  wire \__uuf__._0798_ ;
  wire \__uuf__._0799_ ;
  wire \__uuf__._0800_ ;
  wire \__uuf__._0801_ ;
  wire \__uuf__._0802_ ;
  wire \__uuf__._0803_ ;
  wire \__uuf__._0804_ ;
  wire \__uuf__._0805_ ;
  wire \__uuf__._0806_ ;
  wire \__uuf__._0807_ ;
  wire \__uuf__._0808_ ;
  wire \__uuf__._0809_ ;
  wire \__uuf__._0810_ ;
  wire \__uuf__._0811_ ;
  wire \__uuf__._0812_ ;
  wire \__uuf__._0813_ ;
  wire \__uuf__._0814_ ;
  wire \__uuf__._0815_ ;
  wire \__uuf__._0816_ ;
  wire \__uuf__._0817_ ;
  wire \__uuf__._0818_ ;
  wire \__uuf__._0819_ ;
  wire \__uuf__._0820_ ;
  wire \__uuf__._0821_ ;
  wire \__uuf__._0822_ ;
  wire \__uuf__._0823_ ;
  wire \__uuf__._0824_ ;
  wire \__uuf__._0825_ ;
  wire \__uuf__._0826_ ;
  wire \__uuf__._0827_ ;
  wire \__uuf__._0828_ ;
  wire \__uuf__._0829_ ;
  wire \__uuf__._0830_ ;
  wire \__uuf__._0831_ ;
  wire \__uuf__._0832_ ;
  wire \__uuf__._0833_ ;
  wire \__uuf__._0834_ ;
  wire \__uuf__._0835_ ;
  wire \__uuf__._0836_ ;
  wire \__uuf__._0837_ ;
  wire \__uuf__._0838_ ;
  wire \__uuf__._0839_ ;
  wire \__uuf__._0840_ ;
  wire \__uuf__._0841_ ;
  wire \__uuf__._0842_ ;
  wire \__uuf__._0843_ ;
  wire \__uuf__._0844_ ;
  wire \__uuf__._0845_ ;
  wire \__uuf__._0846_ ;
  wire \__uuf__._0847_ ;
  wire \__uuf__._0848_ ;
  wire \__uuf__._0849_ ;
  wire \__uuf__._0850_ ;
  wire \__uuf__._0851_ ;
  wire \__uuf__._0852_ ;
  wire \__uuf__._0853_ ;
  wire \__uuf__._0854_ ;
  wire \__uuf__._0855_ ;
  wire \__uuf__._0856_ ;
  wire \__uuf__._0857_ ;
  wire \__uuf__._0858_ ;
  wire \__uuf__._0859_ ;
  wire \__uuf__._0860_ ;
  wire \__uuf__._0861_ ;
  wire \__uuf__._0862_ ;
  wire \__uuf__._0863_ ;
  wire \__uuf__._0864_ ;
  wire \__uuf__._0865_ ;
  wire \__uuf__._0866_ ;
  wire \__uuf__._0867_ ;
  wire \__uuf__._0868_ ;
  wire \__uuf__._0869_ ;
  wire \__uuf__._0870_ ;
  wire \__uuf__._0871_ ;
  wire \__uuf__._0872_ ;
  wire \__uuf__._0873_ ;
  wire \__uuf__._0874_ ;
  wire \__uuf__._0875_ ;
  wire \__uuf__._0876_ ;
  wire \__uuf__._0877_ ;
  wire \__uuf__._0878_ ;
  wire \__uuf__._0879_ ;
  wire \__uuf__._0880_ ;
  wire \__uuf__._0881_ ;
  wire \__uuf__.__clk_source__ ;
  wire \__uuf__.count[0] ;
  wire \__uuf__.count[1] ;
  wire \__uuf__.count[2] ;
  wire \__uuf__.count[3] ;
  wire \__uuf__.count[4] ;
  wire \__uuf__.count[5] ;
  wire \__uuf__.fsm.newstate[0] ;
  wire \__uuf__.fsm.newstate[1] ;
  wire \__uuf__.fsm.state[0] ;
  wire \__uuf__.fsm.state[1] ;
  wire \__uuf__.multiplier.csa0.sc ;
  wire \__uuf__.multiplier.csa0.sum ;
  wire \__uuf__.multiplier.csa0.y ;
  wire \__uuf__.multiplier.pp[10] ;
  wire \__uuf__.multiplier.pp[11] ;
  wire \__uuf__.multiplier.pp[12] ;
  wire \__uuf__.multiplier.pp[13] ;
  wire \__uuf__.multiplier.pp[14] ;
  wire \__uuf__.multiplier.pp[15] ;
  wire \__uuf__.multiplier.pp[16] ;
  wire \__uuf__.multiplier.pp[17] ;
  wire \__uuf__.multiplier.pp[18] ;
  wire \__uuf__.multiplier.pp[19] ;
  wire \__uuf__.multiplier.pp[20] ;
  wire \__uuf__.multiplier.pp[21] ;
  wire \__uuf__.multiplier.pp[22] ;
  wire \__uuf__.multiplier.pp[23] ;
  wire \__uuf__.multiplier.pp[24] ;
  wire \__uuf__.multiplier.pp[25] ;
  wire \__uuf__.multiplier.pp[26] ;
  wire \__uuf__.multiplier.pp[27] ;
  wire \__uuf__.multiplier.pp[28] ;
  wire \__uuf__.multiplier.pp[29] ;
  wire \__uuf__.multiplier.pp[2] ;
  wire \__uuf__.multiplier.pp[30] ;
  wire \__uuf__.multiplier.pp[31] ;
  wire \__uuf__.multiplier.pp[3] ;
  wire \__uuf__.multiplier.pp[4] ;
  wire \__uuf__.multiplier.pp[5] ;
  wire \__uuf__.multiplier.pp[6] ;
  wire \__uuf__.multiplier.pp[7] ;
  wire \__uuf__.multiplier.pp[8] ;
  wire \__uuf__.multiplier.pp[9] ;
  wire \__uuf__.multiplier.tcmp.z ;
  wire \__uuf__.multiplier.y ;
  wire \__uuf__.shifter.shiftreg[0] ;
  wire \__uuf__.shifter.shiftreg[10] ;
  wire \__uuf__.shifter.shiftreg[11] ;
  wire \__uuf__.shifter.shiftreg[12] ;
  wire \__uuf__.shifter.shiftreg[13] ;
  wire \__uuf__.shifter.shiftreg[14] ;
  wire \__uuf__.shifter.shiftreg[15] ;
  wire \__uuf__.shifter.shiftreg[16] ;
  wire \__uuf__.shifter.shiftreg[17] ;
  wire \__uuf__.shifter.shiftreg[18] ;
  wire \__uuf__.shifter.shiftreg[19] ;
  wire \__uuf__.shifter.shiftreg[1] ;
  wire \__uuf__.shifter.shiftreg[20] ;
  wire \__uuf__.shifter.shiftreg[21] ;
  wire \__uuf__.shifter.shiftreg[22] ;
  wire \__uuf__.shifter.shiftreg[23] ;
  wire \__uuf__.shifter.shiftreg[24] ;
  wire \__uuf__.shifter.shiftreg[25] ;
  wire \__uuf__.shifter.shiftreg[26] ;
  wire \__uuf__.shifter.shiftreg[27] ;
  wire \__uuf__.shifter.shiftreg[28] ;
  wire \__uuf__.shifter.shiftreg[29] ;
  wire \__uuf__.shifter.shiftreg[2] ;
  wire \__uuf__.shifter.shiftreg[30] ;
  wire \__uuf__.shifter.shiftreg[31] ;
  wire \__uuf__.shifter.shiftreg[32] ;
  wire \__uuf__.shifter.shiftreg[33] ;
  wire \__uuf__.shifter.shiftreg[34] ;
  wire \__uuf__.shifter.shiftreg[35] ;
  wire \__uuf__.shifter.shiftreg[36] ;
  wire \__uuf__.shifter.shiftreg[37] ;
  wire \__uuf__.shifter.shiftreg[38] ;
  wire \__uuf__.shifter.shiftreg[39] ;
  wire \__uuf__.shifter.shiftreg[3] ;
  wire \__uuf__.shifter.shiftreg[40] ;
  wire \__uuf__.shifter.shiftreg[41] ;
  wire \__uuf__.shifter.shiftreg[42] ;
  wire \__uuf__.shifter.shiftreg[43] ;
  wire \__uuf__.shifter.shiftreg[44] ;
  wire \__uuf__.shifter.shiftreg[45] ;
  wire \__uuf__.shifter.shiftreg[46] ;
  wire \__uuf__.shifter.shiftreg[47] ;
  wire \__uuf__.shifter.shiftreg[48] ;
  wire \__uuf__.shifter.shiftreg[49] ;
  wire \__uuf__.shifter.shiftreg[4] ;
  wire \__uuf__.shifter.shiftreg[50] ;
  wire \__uuf__.shifter.shiftreg[51] ;
  wire \__uuf__.shifter.shiftreg[52] ;
  wire \__uuf__.shifter.shiftreg[53] ;
  wire \__uuf__.shifter.shiftreg[54] ;
  wire \__uuf__.shifter.shiftreg[55] ;
  wire \__uuf__.shifter.shiftreg[56] ;
  wire \__uuf__.shifter.shiftreg[57] ;
  wire \__uuf__.shifter.shiftreg[58] ;
  wire \__uuf__.shifter.shiftreg[59] ;
  wire \__uuf__.shifter.shiftreg[5] ;
  wire \__uuf__.shifter.shiftreg[60] ;
  wire \__uuf__.shifter.shiftreg[61] ;
  wire \__uuf__.shifter.shiftreg[62] ;
  wire \__uuf__.shifter.shiftreg[63] ;
  wire \__uuf__.shifter.shiftreg[6] ;
  wire \__uuf__.shifter.shiftreg[7] ;
  wire \__uuf__.shifter.shiftreg[8] ;
  wire \__uuf__.shifter.shiftreg[9] ;
  input clk;
  output done;
  input [31:0] mc;
  input [31:0] mp;
  output [63:0] prod;
  input rst;
  input shift;
  input sin;
  output sout;
  input start;
  input tck;
  input test;

  sky130_fd_sc_hd__and2_4
  _0862_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_5__.sout ),
    .X(_0587_)
  );


  sky130_fd_sc_hd__a21o_4
  _0863_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_6__.dout ),
    .B1(_0587_),
    .X(_0191_)
  );


  sky130_fd_sc_hd__and2_4
  _0864_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_7__.sout ),
    .X(_0588_)
  );


  sky130_fd_sc_hd__a21o_4
  _0865_
  (
    .A1(_0463_),
    .A2(mc[7]),
    .B1(_0588_),
    .X(\__BoundaryScanRegister_input_7__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _0866_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_6__.sout ),
    .X(_0589_)
  );


  sky130_fd_sc_hd__a21o_4
  _0867_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_7__.dout ),
    .B1(_0589_),
    .X(_0192_)
  );


  sky130_fd_sc_hd__and2_4
  _0868_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_8__.sout ),
    .X(_0590_)
  );


  sky130_fd_sc_hd__a21o_4
  _0869_
  (
    .A1(_0463_),
    .A2(mc[8]),
    .B1(_0590_),
    .X(\__BoundaryScanRegister_input_8__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _0870_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_7__.sout ),
    .X(_0591_)
  );


  sky130_fd_sc_hd__a21o_4
  _0871_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_8__.dout ),
    .B1(_0591_),
    .X(_0193_)
  );


  sky130_fd_sc_hd__and2_4
  _0872_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_10__.sin ),
    .X(_0592_)
  );


  sky130_fd_sc_hd__a21o_4
  _0873_
  (
    .A1(_0463_),
    .A2(mc[9]),
    .B1(_0592_),
    .X(\__BoundaryScanRegister_input_9__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _0874_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_8__.sout ),
    .X(_0593_)
  );


  sky130_fd_sc_hd__a21o_4
  _0875_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_9__.dout ),
    .B1(_0593_),
    .X(_0194_)
  );


  sky130_fd_sc_hd__and2_4
  _0876_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_100__.sin ),
    .X(_0594_)
  );


  sky130_fd_sc_hd__a21o_4
  _0877_
  (
    .A1(_0462_),
    .A2(prod[35]),
    .B1(_0594_),
    .X(_0195_)
  );


  sky130_fd_sc_hd__and2_4
  _0878_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_100__.sout ),
    .X(_0595_)
  );


  sky130_fd_sc_hd__a21o_4
  _0879_
  (
    .A1(_0462_),
    .A2(prod[36]),
    .B1(_0595_),
    .X(_0196_)
  );


  sky130_fd_sc_hd__and2_4
  _0880_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_101__.sout ),
    .X(_0596_)
  );


  sky130_fd_sc_hd__a21o_4
  _0881_
  (
    .A1(_0462_),
    .A2(prod[37]),
    .B1(_0596_),
    .X(_0197_)
  );


  sky130_fd_sc_hd__and2_4
  _0882_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_102__.sout ),
    .X(_0597_)
  );


  sky130_fd_sc_hd__a21o_4
  _0883_
  (
    .A1(_0462_),
    .A2(prod[38]),
    .B1(_0597_),
    .X(_0198_)
  );


  sky130_fd_sc_hd__and2_4
  _0884_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_103__.sout ),
    .X(_0598_)
  );


  sky130_fd_sc_hd__a21o_4
  _0885_
  (
    .A1(_0462_),
    .A2(prod[39]),
    .B1(_0598_),
    .X(_0199_)
  );


  sky130_fd_sc_hd__and2_4
  _0886_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_104__.sout ),
    .X(_0599_)
  );


  sky130_fd_sc_hd__a21o_4
  _0887_
  (
    .A1(_0462_),
    .A2(prod[40]),
    .B1(_0599_),
    .X(_0200_)
  );


  sky130_fd_sc_hd__and2_4
  _0888_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_105__.sout ),
    .X(_0600_)
  );


  sky130_fd_sc_hd__a21o_4
  _0889_
  (
    .A1(_0462_),
    .A2(prod[41]),
    .B1(_0600_),
    .X(_0201_)
  );


  sky130_fd_sc_hd__and2_4
  _0890_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_106__.sout ),
    .X(_0601_)
  );


  sky130_fd_sc_hd__a21o_4
  _0891_
  (
    .A1(_0462_),
    .A2(prod[42]),
    .B1(_0601_),
    .X(_0202_)
  );


  sky130_fd_sc_hd__and2_4
  _0892_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_107__.sout ),
    .X(_0602_)
  );


  sky130_fd_sc_hd__a21o_4
  _0893_
  (
    .A1(_0462_),
    .A2(prod[43]),
    .B1(_0602_),
    .X(_0203_)
  );


  sky130_fd_sc_hd__and2_4
  _0894_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_108__.sout ),
    .X(_0603_)
  );


  sky130_fd_sc_hd__a21o_4
  _0895_
  (
    .A1(_0462_),
    .A2(prod[44]),
    .B1(_0603_),
    .X(_0204_)
  );


  sky130_fd_sc_hd__and2_4
  _0896_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_109__.sout ),
    .X(_0604_)
  );


  sky130_fd_sc_hd__a21o_4
  _0897_
  (
    .A1(_0462_),
    .A2(prod[45]),
    .B1(_0604_),
    .X(_0205_)
  );


  sky130_fd_sc_hd__and2_4
  _0898_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_110__.sout ),
    .X(_0605_)
  );


  sky130_fd_sc_hd__a21o_4
  _0899_
  (
    .A1(_0462_),
    .A2(prod[46]),
    .B1(_0605_),
    .X(_0206_)
  );


  sky130_fd_sc_hd__and2_4
  _0900_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_111__.sout ),
    .X(_0606_)
  );


  sky130_fd_sc_hd__a21o_4
  _0901_
  (
    .A1(_0462_),
    .A2(prod[47]),
    .B1(_0606_),
    .X(_0207_)
  );


  sky130_fd_sc_hd__and2_4
  _0902_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_112__.sout ),
    .X(_0607_)
  );


  sky130_fd_sc_hd__a21o_4
  _0903_
  (
    .A1(_0462_),
    .A2(prod[48]),
    .B1(_0607_),
    .X(_0208_)
  );


  sky130_fd_sc_hd__and2_4
  _0904_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_113__.sout ),
    .X(_0608_)
  );


  sky130_fd_sc_hd__a21o_4
  _0905_
  (
    .A1(_0462_),
    .A2(prod[49]),
    .B1(_0608_),
    .X(_0209_)
  );


  sky130_fd_sc_hd__and2_4
  _0906_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_114__.sout ),
    .X(_0609_)
  );


  sky130_fd_sc_hd__a21o_4
  _0907_
  (
    .A1(_0462_),
    .A2(prod[50]),
    .B1(_0609_),
    .X(_0210_)
  );


  sky130_fd_sc_hd__and2_4
  _0908_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_115__.sout ),
    .X(_0610_)
  );


  sky130_fd_sc_hd__a21o_4
  _0909_
  (
    .A1(_0462_),
    .A2(prod[51]),
    .B1(_0610_),
    .X(_0211_)
  );


  sky130_fd_sc_hd__and2_4
  _0910_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_116__.sout ),
    .X(_0611_)
  );


  sky130_fd_sc_hd__a21o_4
  _0911_
  (
    .A1(_0462_),
    .A2(prod[52]),
    .B1(_0611_),
    .X(_0212_)
  );


  sky130_fd_sc_hd__and2_4
  _0912_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_117__.sout ),
    .X(_0612_)
  );


  sky130_fd_sc_hd__a21o_4
  _0913_
  (
    .A1(_0462_),
    .A2(prod[53]),
    .B1(_0612_),
    .X(_0213_)
  );


  sky130_fd_sc_hd__and2_4
  _0914_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_118__.sout ),
    .X(_0613_)
  );


  sky130_fd_sc_hd__a21o_4
  _0915_
  (
    .A1(_0462_),
    .A2(prod[54]),
    .B1(_0613_),
    .X(_0214_)
  );


  sky130_fd_sc_hd__and2_4
  _0916_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_119__.sout ),
    .X(_0614_)
  );


  sky130_fd_sc_hd__a21o_4
  _0917_
  (
    .A1(_0462_),
    .A2(prod[55]),
    .B1(_0614_),
    .X(_0215_)
  );


  sky130_fd_sc_hd__and2_4
  _0918_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_120__.sout ),
    .X(_0615_)
  );


  sky130_fd_sc_hd__a21o_4
  _0919_
  (
    .A1(_0462_),
    .A2(prod[56]),
    .B1(_0615_),
    .X(_0216_)
  );


  sky130_fd_sc_hd__and2_4
  _0920_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_121__.sout ),
    .X(_0616_)
  );


  sky130_fd_sc_hd__a21o_4
  _0921_
  (
    .A1(_0462_),
    .A2(prod[57]),
    .B1(_0616_),
    .X(_0217_)
  );


  sky130_fd_sc_hd__and2_4
  _0922_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_122__.sout ),
    .X(_0617_)
  );


  sky130_fd_sc_hd__a21o_4
  _0923_
  (
    .A1(_0462_),
    .A2(prod[58]),
    .B1(_0617_),
    .X(_0218_)
  );


  sky130_fd_sc_hd__and2_4
  _0924_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_123__.sout ),
    .X(_0618_)
  );


  sky130_fd_sc_hd__a21o_4
  _0925_
  (
    .A1(_0462_),
    .A2(prod[59]),
    .B1(_0618_),
    .X(_0219_)
  );


  sky130_fd_sc_hd__and2_4
  _0926_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_124__.sout ),
    .X(_0619_)
  );


  sky130_fd_sc_hd__a21o_4
  _0927_
  (
    .A1(_0462_),
    .A2(prod[60]),
    .B1(_0619_),
    .X(_0220_)
  );


  sky130_fd_sc_hd__and2_4
  _0928_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_125__.sout ),
    .X(_0620_)
  );


  sky130_fd_sc_hd__a21o_4
  _0929_
  (
    .A1(_0462_),
    .A2(prod[61]),
    .B1(_0620_),
    .X(_0221_)
  );


  sky130_fd_sc_hd__and2_4
  _0930_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_126__.sout ),
    .X(_0621_)
  );


  sky130_fd_sc_hd__a21o_4
  _0931_
  (
    .A1(_0462_),
    .A2(prod[62]),
    .B1(_0621_),
    .X(_0222_)
  );


  sky130_fd_sc_hd__and2_4
  _0932_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_127__.sout ),
    .X(_0622_)
  );


  sky130_fd_sc_hd__a21o_4
  _0933_
  (
    .A1(_0462_),
    .A2(prod[63]),
    .B1(_0622_),
    .X(_0223_)
  );


  sky130_fd_sc_hd__and2_4
  _0934_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_128__.sout ),
    .X(_0623_)
  );


  sky130_fd_sc_hd__a21o_4
  _0935_
  (
    .A1(_0462_),
    .A2(done),
    .B1(_0623_),
    .X(_0224_)
  );


  sky130_fd_sc_hd__and2_4
  _0936_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_65__.sin ),
    .X(_0624_)
  );


  sky130_fd_sc_hd__a21o_4
  _0937_
  (
    .A1(_0462_),
    .A2(prod[0]),
    .B1(_0624_),
    .X(_0225_)
  );


  sky130_fd_sc_hd__and2_4
  _0938_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_65__.sout ),
    .X(_0625_)
  );


  sky130_fd_sc_hd__a21o_4
  _0939_
  (
    .A1(_0462_),
    .A2(prod[1]),
    .B1(_0625_),
    .X(_0226_)
  );


  sky130_fd_sc_hd__and2_4
  _0940_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_66__.sout ),
    .X(_0626_)
  );


  sky130_fd_sc_hd__a21o_4
  _0941_
  (
    .A1(_0462_),
    .A2(prod[2]),
    .B1(_0626_),
    .X(_0227_)
  );


  sky130_fd_sc_hd__and2_4
  _0942_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_67__.sout ),
    .X(_0627_)
  );


  sky130_fd_sc_hd__a21o_4
  _0943_
  (
    .A1(_0462_),
    .A2(prod[3]),
    .B1(_0627_),
    .X(_0228_)
  );


  sky130_fd_sc_hd__and2_4
  _0944_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_68__.sout ),
    .X(_0628_)
  );


  sky130_fd_sc_hd__a21o_4
  _0945_
  (
    .A1(_0462_),
    .A2(prod[4]),
    .B1(_0628_),
    .X(_0229_)
  );


  sky130_fd_sc_hd__and2_4
  _0946_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_69__.sout ),
    .X(_0629_)
  );


  sky130_fd_sc_hd__a21o_4
  _0947_
  (
    .A1(_0462_),
    .A2(prod[5]),
    .B1(_0629_),
    .X(_0230_)
  );


  sky130_fd_sc_hd__and2_4
  _0948_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_70__.sout ),
    .X(_0630_)
  );


  sky130_fd_sc_hd__a21o_4
  _0949_
  (
    .A1(_0462_),
    .A2(prod[6]),
    .B1(_0630_),
    .X(_0231_)
  );


  sky130_fd_sc_hd__and2_4
  _0950_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_71__.sout ),
    .X(_0631_)
  );


  sky130_fd_sc_hd__a21o_4
  _0951_
  (
    .A1(_0462_),
    .A2(prod[7]),
    .B1(_0631_),
    .X(_0232_)
  );


  sky130_fd_sc_hd__and2_4
  _0952_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_72__.sout ),
    .X(_0632_)
  );


  sky130_fd_sc_hd__a21o_4
  _0953_
  (
    .A1(_0462_),
    .A2(prod[8]),
    .B1(_0632_),
    .X(_0233_)
  );


  sky130_fd_sc_hd__and2_4
  _0954_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_73__.sout ),
    .X(_0633_)
  );


  sky130_fd_sc_hd__a21o_4
  _0955_
  (
    .A1(_0462_),
    .A2(prod[9]),
    .B1(_0633_),
    .X(_0234_)
  );


  sky130_fd_sc_hd__and2_4
  _0956_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_74__.sout ),
    .X(_0634_)
  );


  sky130_fd_sc_hd__a21o_4
  _0957_
  (
    .A1(_0462_),
    .A2(prod[10]),
    .B1(_0634_),
    .X(_0235_)
  );


  sky130_fd_sc_hd__and2_4
  _0958_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_75__.sout ),
    .X(_0635_)
  );


  sky130_fd_sc_hd__a21o_4
  _0959_
  (
    .A1(_0462_),
    .A2(prod[11]),
    .B1(_0635_),
    .X(_0236_)
  );


  sky130_fd_sc_hd__and2_4
  _0960_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_76__.sout ),
    .X(_0636_)
  );


  sky130_fd_sc_hd__a21o_4
  _0961_
  (
    .A1(_0462_),
    .A2(prod[12]),
    .B1(_0636_),
    .X(_0237_)
  );


  sky130_fd_sc_hd__and2_4
  _0962_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_77__.sout ),
    .X(_0637_)
  );


  sky130_fd_sc_hd__a21o_4
  _0963_
  (
    .A1(_0462_),
    .A2(prod[13]),
    .B1(_0637_),
    .X(_0238_)
  );


  sky130_fd_sc_hd__and2_4
  _0964_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_78__.sout ),
    .X(_0638_)
  );


  sky130_fd_sc_hd__a21o_4
  _0965_
  (
    .A1(_0462_),
    .A2(prod[14]),
    .B1(_0638_),
    .X(_0239_)
  );


  sky130_fd_sc_hd__and2_4
  _0966_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_79__.sout ),
    .X(_0639_)
  );


  sky130_fd_sc_hd__a21o_4
  _0967_
  (
    .A1(_0462_),
    .A2(prod[15]),
    .B1(_0639_),
    .X(_0240_)
  );


  sky130_fd_sc_hd__and2_4
  _0968_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_80__.sout ),
    .X(_0640_)
  );


  sky130_fd_sc_hd__a21o_4
  _0969_
  (
    .A1(_0462_),
    .A2(prod[16]),
    .B1(_0640_),
    .X(_0241_)
  );


  sky130_fd_sc_hd__and2_4
  _0970_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_81__.sout ),
    .X(_0641_)
  );


  sky130_fd_sc_hd__a21o_4
  _0971_
  (
    .A1(_0462_),
    .A2(prod[17]),
    .B1(_0641_),
    .X(_0242_)
  );


  sky130_fd_sc_hd__and2_4
  _0972_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_82__.sout ),
    .X(_0642_)
  );


  sky130_fd_sc_hd__a21o_4
  _0973_
  (
    .A1(_0462_),
    .A2(prod[18]),
    .B1(_0642_),
    .X(_0243_)
  );


  sky130_fd_sc_hd__and2_4
  _0974_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_83__.sout ),
    .X(_0643_)
  );


  sky130_fd_sc_hd__a21o_4
  _0975_
  (
    .A1(_0462_),
    .A2(prod[19]),
    .B1(_0643_),
    .X(_0244_)
  );


  sky130_fd_sc_hd__and2_4
  _0976_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_84__.sout ),
    .X(_0644_)
  );


  sky130_fd_sc_hd__a21o_4
  _0977_
  (
    .A1(_0462_),
    .A2(prod[20]),
    .B1(_0644_),
    .X(_0245_)
  );


  sky130_fd_sc_hd__and2_4
  _0978_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_85__.sout ),
    .X(_0645_)
  );


  sky130_fd_sc_hd__a21o_4
  _0979_
  (
    .A1(_0462_),
    .A2(prod[21]),
    .B1(_0645_),
    .X(_0246_)
  );


  sky130_fd_sc_hd__and2_4
  _0980_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_86__.sout ),
    .X(_0646_)
  );


  sky130_fd_sc_hd__a21o_4
  _0981_
  (
    .A1(_0462_),
    .A2(prod[22]),
    .B1(_0646_),
    .X(_0247_)
  );


  sky130_fd_sc_hd__and2_4
  _0982_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_87__.sout ),
    .X(_0647_)
  );


  sky130_fd_sc_hd__a21o_4
  _0983_
  (
    .A1(_0462_),
    .A2(prod[23]),
    .B1(_0647_),
    .X(_0248_)
  );


  sky130_fd_sc_hd__and2_4
  _0984_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_88__.sout ),
    .X(_0648_)
  );


  sky130_fd_sc_hd__a21o_4
  _0985_
  (
    .A1(_0462_),
    .A2(prod[24]),
    .B1(_0648_),
    .X(_0249_)
  );


  sky130_fd_sc_hd__and2_4
  _0986_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_89__.sout ),
    .X(_0649_)
  );


  sky130_fd_sc_hd__a21o_4
  _0987_
  (
    .A1(_0462_),
    .A2(prod[25]),
    .B1(_0649_),
    .X(_0250_)
  );


  sky130_fd_sc_hd__and2_4
  _0988_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_90__.sout ),
    .X(_0650_)
  );


  sky130_fd_sc_hd__a21o_4
  _0989_
  (
    .A1(_0462_),
    .A2(prod[26]),
    .B1(_0650_),
    .X(_0251_)
  );


  sky130_fd_sc_hd__and2_4
  _0990_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_91__.sout ),
    .X(_0651_)
  );


  sky130_fd_sc_hd__a21o_4
  _0991_
  (
    .A1(_0462_),
    .A2(prod[27]),
    .B1(_0651_),
    .X(_0252_)
  );


  sky130_fd_sc_hd__and2_4
  _0992_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_92__.sout ),
    .X(_0652_)
  );


  sky130_fd_sc_hd__a21o_4
  _0993_
  (
    .A1(_0462_),
    .A2(prod[28]),
    .B1(_0652_),
    .X(_0253_)
  );


  sky130_fd_sc_hd__and2_4
  _0994_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_93__.sout ),
    .X(_0653_)
  );


  sky130_fd_sc_hd__a21o_4
  _0995_
  (
    .A1(_0462_),
    .A2(prod[29]),
    .B1(_0653_),
    .X(_0254_)
  );


  sky130_fd_sc_hd__and2_4
  _0996_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_94__.sout ),
    .X(_0654_)
  );


  sky130_fd_sc_hd__a21o_4
  _0997_
  (
    .A1(_0462_),
    .A2(prod[30]),
    .B1(_0654_),
    .X(_0255_)
  );


  sky130_fd_sc_hd__and2_4
  _0998_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_95__.sout ),
    .X(_0655_)
  );


  sky130_fd_sc_hd__a21o_4
  _0999_
  (
    .A1(_0462_),
    .A2(prod[31]),
    .B1(_0655_),
    .X(_0256_)
  );


  sky130_fd_sc_hd__and2_4
  _1000_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_96__.sout ),
    .X(_0656_)
  );


  sky130_fd_sc_hd__a21o_4
  _1001_
  (
    .A1(_0462_),
    .A2(prod[32]),
    .B1(_0656_),
    .X(_0257_)
  );


  sky130_fd_sc_hd__and2_4
  _1002_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_97__.sout ),
    .X(_0657_)
  );


  sky130_fd_sc_hd__a21o_4
  _1003_
  (
    .A1(_0462_),
    .A2(prod[33]),
    .B1(_0657_),
    .X(_0258_)
  );


  sky130_fd_sc_hd__and2_4
  _1004_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_output_98__.sout ),
    .X(_0658_)
  );


  sky130_fd_sc_hd__a21o_4
  _1005_
  (
    .A1(_0462_),
    .A2(prod[34]),
    .B1(_0658_),
    .X(_0259_)
  );


  sky130_fd_sc_hd__and2_4
  _1006_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_64__.sout ),
    .X(_0659_)
  );


  sky130_fd_sc_hd__a21o_4
  _1007_
  (
    .A1(_0462_),
    .A2(\__uuf__._0095_ ),
    .B1(_0659_),
    .X(_0342_)
  );


  sky130_fd_sc_hd__and2_4
  _1008_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[0] ),
    .X(_0660_)
  );


  sky130_fd_sc_hd__a21o_4
  _1009_
  (
    .A1(_0462_),
    .A2(\__uuf__._0106_ ),
    .B1(_0660_),
    .X(_0343_)
  );


  sky130_fd_sc_hd__and2_4
  _1010_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[1] ),
    .X(_0661_)
  );


  sky130_fd_sc_hd__a21o_4
  _1011_
  (
    .A1(_0462_),
    .A2(\__uuf__._0117_ ),
    .B1(_0661_),
    .X(_0344_)
  );


  sky130_fd_sc_hd__and2_4
  _1012_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[2] ),
    .X(_0662_)
  );


  sky130_fd_sc_hd__a21o_4
  _1013_
  (
    .A1(_0462_),
    .A2(\__uuf__._0128_ ),
    .B1(_0662_),
    .X(_0345_)
  );


  sky130_fd_sc_hd__and2_4
  _1014_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[3] ),
    .X(_0663_)
  );


  sky130_fd_sc_hd__a21o_4
  _1015_
  (
    .A1(_0462_),
    .A2(\__uuf__._0139_ ),
    .B1(_0663_),
    .X(_0346_)
  );


  sky130_fd_sc_hd__and2_4
  _1016_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[4] ),
    .X(_0664_)
  );


  sky130_fd_sc_hd__a21o_4
  _1017_
  (
    .A1(_0462_),
    .A2(\__uuf__._0150_ ),
    .B1(_0664_),
    .X(_0347_)
  );


  sky130_fd_sc_hd__and2_4
  _1018_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[5] ),
    .X(_0665_)
  );


  sky130_fd_sc_hd__a21o_4
  _1019_
  (
    .A1(_0462_),
    .A2(\__uuf__._0155_ ),
    .B1(_0665_),
    .X(_0348_)
  );


  sky130_fd_sc_hd__and2_4
  _1020_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[6] ),
    .X(_0666_)
  );


  sky130_fd_sc_hd__a21o_4
  _1021_
  (
    .A1(_0462_),
    .A2(\__uuf__._0156_ ),
    .B1(_0666_),
    .X(_0349_)
  );


  sky130_fd_sc_hd__and2_4
  _1022_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[7] ),
    .X(_0667_)
  );


  sky130_fd_sc_hd__a21o_4
  _1023_
  (
    .A1(_0462_),
    .A2(\__uuf__._0157_ ),
    .B1(_0667_),
    .X(_0350_)
  );


  sky130_fd_sc_hd__and2_4
  _1024_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[8] ),
    .X(_0668_)
  );


  sky130_fd_sc_hd__a21o_4
  _1025_
  (
    .A1(_0462_),
    .A2(\__uuf__._0158_ ),
    .B1(_0668_),
    .X(_0351_)
  );


  sky130_fd_sc_hd__and2_4
  _1026_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[9] ),
    .X(_0669_)
  );


  sky130_fd_sc_hd__a21o_4
  _1027_
  (
    .A1(_0462_),
    .A2(\__uuf__._0096_ ),
    .B1(_0669_),
    .X(_0352_)
  );


  sky130_fd_sc_hd__and2_4
  _1028_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[10] ),
    .X(_0670_)
  );


  sky130_fd_sc_hd__a21o_4
  _1029_
  (
    .A1(_0462_),
    .A2(\__uuf__._0097_ ),
    .B1(_0670_),
    .X(_0353_)
  );


  sky130_fd_sc_hd__and2_4
  _1030_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[11] ),
    .X(_0671_)
  );


  sky130_fd_sc_hd__a21o_4
  _1031_
  (
    .A1(_0462_),
    .A2(\__uuf__._0098_ ),
    .B1(_0671_),
    .X(_0354_)
  );


  sky130_fd_sc_hd__and2_4
  _1032_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[12] ),
    .X(_0672_)
  );


  sky130_fd_sc_hd__a21o_4
  _1033_
  (
    .A1(_0462_),
    .A2(\__uuf__._0099_ ),
    .B1(_0672_),
    .X(_0355_)
  );


  sky130_fd_sc_hd__and2_4
  _1034_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[13] ),
    .X(_0673_)
  );


  sky130_fd_sc_hd__a21o_4
  _1035_
  (
    .A1(_0462_),
    .A2(\__uuf__._0100_ ),
    .B1(_0673_),
    .X(_0356_)
  );


  sky130_fd_sc_hd__and2_4
  _1036_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[14] ),
    .X(_0674_)
  );


  sky130_fd_sc_hd__a21o_4
  _1037_
  (
    .A1(_0462_),
    .A2(\__uuf__._0101_ ),
    .B1(_0674_),
    .X(_0357_)
  );


  sky130_fd_sc_hd__and2_4
  _1038_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[15] ),
    .X(_0675_)
  );


  sky130_fd_sc_hd__a21o_4
  _1039_
  (
    .A1(_0462_),
    .A2(\__uuf__._0102_ ),
    .B1(_0675_),
    .X(_0358_)
  );


  sky130_fd_sc_hd__and2_4
  _1040_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[16] ),
    .X(_0676_)
  );


  sky130_fd_sc_hd__a21o_4
  _1041_
  (
    .A1(_0462_),
    .A2(\__uuf__._0103_ ),
    .B1(_0676_),
    .X(_0359_)
  );


  sky130_fd_sc_hd__and2_4
  _1042_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[17] ),
    .X(_0677_)
  );


  sky130_fd_sc_hd__a21o_4
  _1043_
  (
    .A1(_0462_),
    .A2(\__uuf__._0104_ ),
    .B1(_0677_),
    .X(_0360_)
  );


  sky130_fd_sc_hd__and2_4
  _1044_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[18] ),
    .X(_0678_)
  );


  sky130_fd_sc_hd__a21o_4
  _1045_
  (
    .A1(_0462_),
    .A2(\__uuf__._0105_ ),
    .B1(_0678_),
    .X(_0361_)
  );


  sky130_fd_sc_hd__and2_4
  _1046_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[19] ),
    .X(_0679_)
  );


  sky130_fd_sc_hd__a21o_4
  _1047_
  (
    .A1(_0462_),
    .A2(\__uuf__._0107_ ),
    .B1(_0679_),
    .X(_0362_)
  );


  sky130_fd_sc_hd__and2_4
  _1048_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[20] ),
    .X(_0680_)
  );


  sky130_fd_sc_hd__a21o_4
  _1049_
  (
    .A1(_0462_),
    .A2(\__uuf__._0108_ ),
    .B1(_0680_),
    .X(_0363_)
  );


  sky130_fd_sc_hd__and2_4
  _1050_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[21] ),
    .X(_0681_)
  );


  sky130_fd_sc_hd__a21o_4
  _1051_
  (
    .A1(_0462_),
    .A2(\__uuf__._0109_ ),
    .B1(_0681_),
    .X(_0364_)
  );


  sky130_fd_sc_hd__and2_4
  _1052_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[22] ),
    .X(_0682_)
  );


  sky130_fd_sc_hd__a21o_4
  _1053_
  (
    .A1(_0462_),
    .A2(\__uuf__._0110_ ),
    .B1(_0682_),
    .X(_0365_)
  );


  sky130_fd_sc_hd__and2_4
  _1054_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[23] ),
    .X(_0683_)
  );


  sky130_fd_sc_hd__a21o_4
  _1055_
  (
    .A1(_0462_),
    .A2(\__uuf__._0111_ ),
    .B1(_0683_),
    .X(_0366_)
  );


  sky130_fd_sc_hd__and2_4
  _1056_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[24] ),
    .X(_0684_)
  );


  sky130_fd_sc_hd__a21o_4
  _1057_
  (
    .A1(_0462_),
    .A2(\__uuf__._0112_ ),
    .B1(_0684_),
    .X(_0367_)
  );


  sky130_fd_sc_hd__and2_4
  _1058_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[25] ),
    .X(_0685_)
  );


  sky130_fd_sc_hd__a21o_4
  _1059_
  (
    .A1(_0462_),
    .A2(\__uuf__._0113_ ),
    .B1(_0685_),
    .X(_0368_)
  );


  sky130_fd_sc_hd__and2_4
  _1060_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[26] ),
    .X(_0686_)
  );


  sky130_fd_sc_hd__a21o_4
  _1061_
  (
    .A1(_0462_),
    .A2(\__uuf__._0114_ ),
    .B1(_0686_),
    .X(_0369_)
  );


  sky130_fd_sc_hd__and2_4
  _1062_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[27] ),
    .X(_0687_)
  );


  sky130_fd_sc_hd__a21o_4
  _1063_
  (
    .A1(_0462_),
    .A2(\__uuf__._0115_ ),
    .B1(_0687_),
    .X(_0370_)
  );


  sky130_fd_sc_hd__and2_4
  _1064_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[28] ),
    .X(_0688_)
  );


  sky130_fd_sc_hd__a21o_4
  _1065_
  (
    .A1(_0462_),
    .A2(\__uuf__._0116_ ),
    .B1(_0688_),
    .X(_0371_)
  );


  sky130_fd_sc_hd__and2_4
  _1066_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[29] ),
    .X(_0689_)
  );


  sky130_fd_sc_hd__a21o_4
  _1067_
  (
    .A1(_0462_),
    .A2(\__uuf__._0118_ ),
    .B1(_0689_),
    .X(_0372_)
  );


  sky130_fd_sc_hd__and2_4
  _1068_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[30] ),
    .X(_0690_)
  );


  sky130_fd_sc_hd__a21o_4
  _1069_
  (
    .A1(_0462_),
    .A2(\__uuf__._0119_ ),
    .B1(_0690_),
    .X(_0373_)
  );


  sky130_fd_sc_hd__and2_4
  _1070_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[31] ),
    .X(_0691_)
  );


  sky130_fd_sc_hd__a21o_4
  _1071_
  (
    .A1(_0462_),
    .A2(\__uuf__._0120_ ),
    .B1(_0691_),
    .X(_0374_)
  );


  sky130_fd_sc_hd__and2_4
  _1072_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[32] ),
    .X(_0692_)
  );


  sky130_fd_sc_hd__a21o_4
  _1073_
  (
    .A1(_0462_),
    .A2(\__uuf__._0121_ ),
    .B1(_0692_),
    .X(_0375_)
  );


  sky130_fd_sc_hd__and2_4
  _1074_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[33] ),
    .X(_0693_)
  );


  sky130_fd_sc_hd__a21o_4
  _1075_
  (
    .A1(_0462_),
    .A2(\__uuf__._0122_ ),
    .B1(_0693_),
    .X(_0376_)
  );


  sky130_fd_sc_hd__and2_4
  _1076_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[34] ),
    .X(_0694_)
  );


  sky130_fd_sc_hd__a21o_4
  _1077_
  (
    .A1(_0462_),
    .A2(\__uuf__._0123_ ),
    .B1(_0694_),
    .X(_0377_)
  );


  sky130_fd_sc_hd__and2_4
  _1078_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[35] ),
    .X(_0695_)
  );


  sky130_fd_sc_hd__a21o_4
  _1079_
  (
    .A1(_0462_),
    .A2(\__uuf__._0124_ ),
    .B1(_0695_),
    .X(_0378_)
  );


  sky130_fd_sc_hd__and2_4
  _1080_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[36] ),
    .X(_0696_)
  );


  sky130_fd_sc_hd__a21o_4
  _1081_
  (
    .A1(_0462_),
    .A2(\__uuf__._0125_ ),
    .B1(_0696_),
    .X(_0379_)
  );


  sky130_fd_sc_hd__and2_4
  _1082_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[37] ),
    .X(_0697_)
  );


  sky130_fd_sc_hd__a21o_4
  _1083_
  (
    .A1(_0462_),
    .A2(\__uuf__._0126_ ),
    .B1(_0697_),
    .X(_0380_)
  );


  sky130_fd_sc_hd__and2_4
  _1084_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[38] ),
    .X(_0698_)
  );


  sky130_fd_sc_hd__a21o_4
  _1085_
  (
    .A1(_0462_),
    .A2(\__uuf__._0127_ ),
    .B1(_0698_),
    .X(_0381_)
  );


  sky130_fd_sc_hd__and2_4
  _1086_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[39] ),
    .X(_0699_)
  );


  sky130_fd_sc_hd__a21o_4
  _1087_
  (
    .A1(_0462_),
    .A2(\__uuf__._0129_ ),
    .B1(_0699_),
    .X(_0382_)
  );


  sky130_fd_sc_hd__and2_4
  _1088_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[40] ),
    .X(_0700_)
  );


  sky130_fd_sc_hd__a21o_4
  _1089_
  (
    .A1(_0462_),
    .A2(\__uuf__._0130_ ),
    .B1(_0700_),
    .X(_0383_)
  );


  sky130_fd_sc_hd__and2_4
  _1090_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[41] ),
    .X(_0701_)
  );


  sky130_fd_sc_hd__a21o_4
  _1091_
  (
    .A1(_0462_),
    .A2(\__uuf__._0131_ ),
    .B1(_0701_),
    .X(_0384_)
  );


  sky130_fd_sc_hd__and2_4
  _1092_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[42] ),
    .X(_0702_)
  );


  sky130_fd_sc_hd__a21o_4
  _1093_
  (
    .A1(_0462_),
    .A2(\__uuf__._0132_ ),
    .B1(_0702_),
    .X(_0385_)
  );


  sky130_fd_sc_hd__and2_4
  _1094_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[43] ),
    .X(_0703_)
  );


  sky130_fd_sc_hd__a21o_4
  _1095_
  (
    .A1(_0462_),
    .A2(\__uuf__._0133_ ),
    .B1(_0703_),
    .X(_0386_)
  );


  sky130_fd_sc_hd__and2_4
  _1096_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[44] ),
    .X(_0704_)
  );


  sky130_fd_sc_hd__a21o_4
  _1097_
  (
    .A1(_0462_),
    .A2(\__uuf__._0134_ ),
    .B1(_0704_),
    .X(_0387_)
  );


  sky130_fd_sc_hd__and2_4
  _1098_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[45] ),
    .X(_0705_)
  );


  sky130_fd_sc_hd__a21o_4
  _1099_
  (
    .A1(_0462_),
    .A2(\__uuf__._0135_ ),
    .B1(_0705_),
    .X(_0388_)
  );


  sky130_fd_sc_hd__and2_4
  _1100_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[46] ),
    .X(_0706_)
  );


  sky130_fd_sc_hd__a21o_4
  _1101_
  (
    .A1(_0462_),
    .A2(\__uuf__._0136_ ),
    .B1(_0706_),
    .X(_0389_)
  );


  sky130_fd_sc_hd__and2_4
  _1102_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[47] ),
    .X(_0707_)
  );


  sky130_fd_sc_hd__a21o_4
  _1103_
  (
    .A1(_0462_),
    .A2(\__uuf__._0137_ ),
    .B1(_0707_),
    .X(_0390_)
  );


  sky130_fd_sc_hd__and2_4
  _1104_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[48] ),
    .X(_0708_)
  );


  sky130_fd_sc_hd__a21o_4
  _1105_
  (
    .A1(_0462_),
    .A2(\__uuf__._0138_ ),
    .B1(_0708_),
    .X(_0391_)
  );


  sky130_fd_sc_hd__and2_4
  _1106_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[49] ),
    .X(_0709_)
  );


  sky130_fd_sc_hd__a21o_4
  _1107_
  (
    .A1(_0462_),
    .A2(\__uuf__._0140_ ),
    .B1(_0709_),
    .X(_0392_)
  );


  sky130_fd_sc_hd__and2_4
  _1108_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[50] ),
    .X(_0710_)
  );


  sky130_fd_sc_hd__a21o_4
  _1109_
  (
    .A1(_0462_),
    .A2(\__uuf__._0141_ ),
    .B1(_0710_),
    .X(_0393_)
  );


  sky130_fd_sc_hd__and2_4
  _1110_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[51] ),
    .X(_0711_)
  );


  sky130_fd_sc_hd__a21o_4
  _1111_
  (
    .A1(_0462_),
    .A2(\__uuf__._0142_ ),
    .B1(_0711_),
    .X(_0394_)
  );


  sky130_fd_sc_hd__and2_4
  _1112_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[52] ),
    .X(_0712_)
  );


  sky130_fd_sc_hd__a21o_4
  _1113_
  (
    .A1(_0462_),
    .A2(\__uuf__._0143_ ),
    .B1(_0712_),
    .X(_0395_)
  );


  sky130_fd_sc_hd__and2_4
  _1114_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[53] ),
    .X(_0713_)
  );


  sky130_fd_sc_hd__a21o_4
  _1115_
  (
    .A1(_0462_),
    .A2(\__uuf__._0144_ ),
    .B1(_0713_),
    .X(_0396_)
  );


  sky130_fd_sc_hd__and2_4
  _1116_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[54] ),
    .X(_0714_)
  );


  sky130_fd_sc_hd__a21o_4
  _1117_
  (
    .A1(_0462_),
    .A2(\__uuf__._0145_ ),
    .B1(_0714_),
    .X(_0397_)
  );


  sky130_fd_sc_hd__and2_4
  _1118_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[55] ),
    .X(_0715_)
  );


  sky130_fd_sc_hd__a21o_4
  _1119_
  (
    .A1(_0462_),
    .A2(\__uuf__._0146_ ),
    .B1(_0715_),
    .X(_0398_)
  );


  sky130_fd_sc_hd__and2_4
  _1120_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[56] ),
    .X(_0716_)
  );


  sky130_fd_sc_hd__a21o_4
  _1121_
  (
    .A1(_0462_),
    .A2(\__uuf__._0147_ ),
    .B1(_0716_),
    .X(_0399_)
  );


  sky130_fd_sc_hd__and2_4
  _1122_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[57] ),
    .X(_0717_)
  );


  sky130_fd_sc_hd__a21o_4
  _1123_
  (
    .A1(_0462_),
    .A2(\__uuf__._0148_ ),
    .B1(_0717_),
    .X(_0400_)
  );


  sky130_fd_sc_hd__and2_4
  _1124_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[58] ),
    .X(_0718_)
  );


  sky130_fd_sc_hd__a21o_4
  _1125_
  (
    .A1(_0462_),
    .A2(\__uuf__._0149_ ),
    .B1(_0718_),
    .X(_0401_)
  );


  sky130_fd_sc_hd__and2_4
  _1126_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[59] ),
    .X(_0719_)
  );


  sky130_fd_sc_hd__a21o_4
  _1127_
  (
    .A1(_0462_),
    .A2(\__uuf__._0151_ ),
    .B1(_0719_),
    .X(_0402_)
  );


  sky130_fd_sc_hd__and2_4
  _1128_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[60] ),
    .X(_0720_)
  );


  sky130_fd_sc_hd__a21o_4
  _1129_
  (
    .A1(_0462_),
    .A2(\__uuf__._0152_ ),
    .B1(_0720_),
    .X(_0403_)
  );


  sky130_fd_sc_hd__and2_4
  _1130_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[61] ),
    .X(_0721_)
  );


  sky130_fd_sc_hd__a21o_4
  _1131_
  (
    .A1(_0462_),
    .A2(\__uuf__._0153_ ),
    .B1(_0721_),
    .X(_0404_)
  );


  sky130_fd_sc_hd__and2_4
  _1132_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[62] ),
    .X(_0722_)
  );


  sky130_fd_sc_hd__a21o_4
  _1133_
  (
    .A1(_0462_),
    .A2(\__uuf__._0154_ ),
    .B1(_0722_),
    .X(_0405_)
  );


  sky130_fd_sc_hd__and2_4
  _1134_
  (
    .A(shift),
    .B(\__uuf__.shifter.shiftreg[63] ),
    .X(_0723_)
  );


  sky130_fd_sc_hd__a21o_4
  _1135_
  (
    .A1(_0462_),
    .A2(\__uuf__._0094_ ),
    .B1(_0723_),
    .X(_0406_)
  );


  sky130_fd_sc_hd__and2_4
  _1136_
  (
    .A(shift),
    .B(\__uuf__.multiplier.y ),
    .X(_0724_)
  );


  sky130_fd_sc_hd__a21o_4
  _1137_
  (
    .A1(_0462_),
    .A2(\__uuf__._0082_ ),
    .B1(_0724_),
    .X(_0407_)
  );


  sky130_fd_sc_hd__and2_4
  _1138_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[30] ),
    .X(_0725_)
  );


  sky130_fd_sc_hd__a21o_4
  _1139_
  (
    .A1(_0462_),
    .A2(\__uuf__._0081_ ),
    .B1(_0725_),
    .X(_0408_)
  );


  sky130_fd_sc_hd__and2_4
  _1140_
  (
    .A(shift),
    .B(\__uuf__._0083_ ),
    .X(_0726_)
  );


  sky130_fd_sc_hd__a21o_4
  _1141_
  (
    .A1(_0462_),
    .A2(\__uuf__._0079_ ),
    .B1(_0726_),
    .X(_0409_)
  );


  sky130_fd_sc_hd__and2_4
  _1142_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[29] ),
    .X(_0727_)
  );


  sky130_fd_sc_hd__a21o_4
  _1143_
  (
    .A1(_0462_),
    .A2(\__uuf__._0078_ ),
    .B1(_0727_),
    .X(_0410_)
  );


  sky130_fd_sc_hd__and2_4
  _1144_
  (
    .A(shift),
    .B(\__uuf__._0080_ ),
    .X(_0728_)
  );


  sky130_fd_sc_hd__a21o_4
  _1145_
  (
    .A1(_0462_),
    .A2(\__uuf__._0076_ ),
    .B1(_0728_),
    .X(_0411_)
  );


  sky130_fd_sc_hd__and2_4
  _1146_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[28] ),
    .X(_0729_)
  );


  sky130_fd_sc_hd__a21o_4
  _1147_
  (
    .A1(_0462_),
    .A2(\__uuf__._0075_ ),
    .B1(_0729_),
    .X(_0412_)
  );


  sky130_fd_sc_hd__and2_4
  _1148_
  (
    .A(shift),
    .B(\__uuf__._0077_ ),
    .X(_0730_)
  );


  sky130_fd_sc_hd__a21o_4
  _1149_
  (
    .A1(_0462_),
    .A2(\__uuf__._0073_ ),
    .B1(_0730_),
    .X(_0413_)
  );


  sky130_fd_sc_hd__and2_4
  _1150_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[27] ),
    .X(_0731_)
  );


  sky130_fd_sc_hd__a21o_4
  _1151_
  (
    .A1(_0462_),
    .A2(\__uuf__._0072_ ),
    .B1(_0731_),
    .X(_0414_)
  );


  sky130_fd_sc_hd__and2_4
  _1152_
  (
    .A(shift),
    .B(\__uuf__._0074_ ),
    .X(_0732_)
  );


  sky130_fd_sc_hd__a21o_4
  _1153_
  (
    .A1(_0462_),
    .A2(\__uuf__._0070_ ),
    .B1(_0732_),
    .X(_0415_)
  );


  sky130_fd_sc_hd__and2_4
  _1154_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[26] ),
    .X(_0733_)
  );


  sky130_fd_sc_hd__a21o_4
  _1155_
  (
    .A1(_0462_),
    .A2(\__uuf__._0069_ ),
    .B1(_0733_),
    .X(_0416_)
  );


  sky130_fd_sc_hd__and2_4
  _1156_
  (
    .A(shift),
    .B(\__uuf__._0071_ ),
    .X(_0734_)
  );


  sky130_fd_sc_hd__a21o_4
  _1157_
  (
    .A1(_0462_),
    .A2(\__uuf__._0067_ ),
    .B1(_0734_),
    .X(_0417_)
  );


  sky130_fd_sc_hd__and2_4
  _1158_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[25] ),
    .X(_0735_)
  );


  sky130_fd_sc_hd__a21o_4
  _1159_
  (
    .A1(_0462_),
    .A2(\__uuf__._0066_ ),
    .B1(_0735_),
    .X(_0418_)
  );


  sky130_fd_sc_hd__and2_4
  _1160_
  (
    .A(shift),
    .B(\__uuf__._0068_ ),
    .X(_0736_)
  );


  sky130_fd_sc_hd__a21o_4
  _1161_
  (
    .A1(_0462_),
    .A2(\__uuf__._0064_ ),
    .B1(_0736_),
    .X(_0419_)
  );


  sky130_fd_sc_hd__and2_4
  _1162_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[24] ),
    .X(_0737_)
  );


  sky130_fd_sc_hd__a21o_4
  _1163_
  (
    .A1(_0462_),
    .A2(\__uuf__._0063_ ),
    .B1(_0737_),
    .X(_0420_)
  );


  sky130_fd_sc_hd__and2_4
  _1164_
  (
    .A(shift),
    .B(\__uuf__._0065_ ),
    .X(_0738_)
  );


  sky130_fd_sc_hd__a21o_4
  _1165_
  (
    .A1(_0462_),
    .A2(\__uuf__._0061_ ),
    .B1(_0738_),
    .X(_0421_)
  );


  sky130_fd_sc_hd__and2_4
  _1166_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[23] ),
    .X(_0739_)
  );


  sky130_fd_sc_hd__a21o_4
  _1167_
  (
    .A1(_0462_),
    .A2(\__uuf__._0060_ ),
    .B1(_0739_),
    .X(_0422_)
  );


  sky130_fd_sc_hd__and2_4
  _1168_
  (
    .A(shift),
    .B(\__uuf__._0062_ ),
    .X(_0740_)
  );


  sky130_fd_sc_hd__a21o_4
  _1169_
  (
    .A1(_0462_),
    .A2(\__uuf__._0058_ ),
    .B1(_0740_),
    .X(_0423_)
  );


  sky130_fd_sc_hd__and2_4
  _1170_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[22] ),
    .X(_0741_)
  );


  sky130_fd_sc_hd__a21o_4
  _1171_
  (
    .A1(_0462_),
    .A2(\__uuf__._0057_ ),
    .B1(_0741_),
    .X(_0424_)
  );


  sky130_fd_sc_hd__and2_4
  _1172_
  (
    .A(shift),
    .B(\__uuf__._0059_ ),
    .X(_0742_)
  );


  sky130_fd_sc_hd__a21o_4
  _1173_
  (
    .A1(_0462_),
    .A2(\__uuf__._0055_ ),
    .B1(_0742_),
    .X(_0425_)
  );


  sky130_fd_sc_hd__and2_4
  _1174_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[21] ),
    .X(_0743_)
  );


  sky130_fd_sc_hd__a21o_4
  _1175_
  (
    .A1(_0462_),
    .A2(\__uuf__._0054_ ),
    .B1(_0743_),
    .X(_0426_)
  );


  sky130_fd_sc_hd__and2_4
  _1176_
  (
    .A(shift),
    .B(\__uuf__._0056_ ),
    .X(_0744_)
  );


  sky130_fd_sc_hd__a21o_4
  _1177_
  (
    .A1(_0462_),
    .A2(\__uuf__._0052_ ),
    .B1(_0744_),
    .X(_0427_)
  );


  sky130_fd_sc_hd__and2_4
  _1178_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[20] ),
    .X(_0745_)
  );


  sky130_fd_sc_hd__a21o_4
  _1179_
  (
    .A1(_0462_),
    .A2(\__uuf__._0051_ ),
    .B1(_0745_),
    .X(_0428_)
  );


  sky130_fd_sc_hd__and2_4
  _1180_
  (
    .A(shift),
    .B(\__uuf__._0053_ ),
    .X(_0746_)
  );


  sky130_fd_sc_hd__a21o_4
  _1181_
  (
    .A1(_0462_),
    .A2(\__uuf__._0049_ ),
    .B1(_0746_),
    .X(_0429_)
  );


  sky130_fd_sc_hd__and2_4
  _1182_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[19] ),
    .X(_0747_)
  );


  sky130_fd_sc_hd__a21o_4
  _1183_
  (
    .A1(_0462_),
    .A2(\__uuf__._0048_ ),
    .B1(_0747_),
    .X(_0430_)
  );


  sky130_fd_sc_hd__and2_4
  _1184_
  (
    .A(shift),
    .B(\__uuf__._0050_ ),
    .X(_0748_)
  );


  sky130_fd_sc_hd__a21o_4
  _1185_
  (
    .A1(_0462_),
    .A2(\__uuf__._0046_ ),
    .B1(_0748_),
    .X(_0431_)
  );


  sky130_fd_sc_hd__and2_4
  _1186_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[18] ),
    .X(_0749_)
  );


  sky130_fd_sc_hd__a21o_4
  _1187_
  (
    .A1(_0462_),
    .A2(\__uuf__._0045_ ),
    .B1(_0749_),
    .X(_0432_)
  );


  sky130_fd_sc_hd__and2_4
  _1188_
  (
    .A(shift),
    .B(\__uuf__._0047_ ),
    .X(_0750_)
  );


  sky130_fd_sc_hd__a21o_4
  _1189_
  (
    .A1(_0462_),
    .A2(\__uuf__._0043_ ),
    .B1(_0750_),
    .X(_0433_)
  );


  sky130_fd_sc_hd__and2_4
  _1190_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[17] ),
    .X(_0751_)
  );


  sky130_fd_sc_hd__a21o_4
  _1191_
  (
    .A1(_0462_),
    .A2(\__uuf__._0042_ ),
    .B1(_0751_),
    .X(_0434_)
  );


  sky130_fd_sc_hd__and2_4
  _1192_
  (
    .A(shift),
    .B(\__uuf__._0044_ ),
    .X(_0752_)
  );


  sky130_fd_sc_hd__a21o_4
  _1193_
  (
    .A1(_0462_),
    .A2(\__uuf__._0040_ ),
    .B1(_0752_),
    .X(_0435_)
  );


  sky130_fd_sc_hd__and2_4
  _1194_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[16] ),
    .X(_0753_)
  );


  sky130_fd_sc_hd__a21o_4
  _1195_
  (
    .A1(_0462_),
    .A2(\__uuf__._0039_ ),
    .B1(_0753_),
    .X(_0436_)
  );


  sky130_fd_sc_hd__and2_4
  _1196_
  (
    .A(shift),
    .B(\__uuf__._0041_ ),
    .X(_0754_)
  );


  sky130_fd_sc_hd__a21o_4
  _1197_
  (
    .A1(_0462_),
    .A2(\__uuf__._0037_ ),
    .B1(_0754_),
    .X(_0437_)
  );


  sky130_fd_sc_hd__and2_4
  _1198_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[15] ),
    .X(_0755_)
  );


  sky130_fd_sc_hd__a21o_4
  _1199_
  (
    .A1(_0462_),
    .A2(\__uuf__._0036_ ),
    .B1(_0755_),
    .X(_0438_)
  );


  sky130_fd_sc_hd__and2_4
  _1200_
  (
    .A(shift),
    .B(\__uuf__._0038_ ),
    .X(_0756_)
  );


  sky130_fd_sc_hd__a21o_4
  _1201_
  (
    .A1(_0462_),
    .A2(\__uuf__._0034_ ),
    .B1(_0756_),
    .X(_0439_)
  );


  sky130_fd_sc_hd__and2_4
  _1202_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[14] ),
    .X(_0757_)
  );


  sky130_fd_sc_hd__a21o_4
  _1203_
  (
    .A1(_0462_),
    .A2(\__uuf__._0033_ ),
    .B1(_0757_),
    .X(_0440_)
  );


  sky130_fd_sc_hd__and2_4
  _1204_
  (
    .A(shift),
    .B(\__uuf__._0035_ ),
    .X(_0758_)
  );


  sky130_fd_sc_hd__a21o_4
  _1205_
  (
    .A1(_0462_),
    .A2(\__uuf__._0031_ ),
    .B1(_0758_),
    .X(_0441_)
  );


  sky130_fd_sc_hd__and2_4
  _1206_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[13] ),
    .X(_0759_)
  );


  sky130_fd_sc_hd__a21o_4
  _1207_
  (
    .A1(_0462_),
    .A2(\__uuf__._0030_ ),
    .B1(_0759_),
    .X(_0442_)
  );


  sky130_fd_sc_hd__and2_4
  _1208_
  (
    .A(shift),
    .B(\__uuf__._0032_ ),
    .X(_0760_)
  );


  sky130_fd_sc_hd__a21o_4
  _1209_
  (
    .A1(_0462_),
    .A2(\__uuf__._0028_ ),
    .B1(_0760_),
    .X(_0443_)
  );


  sky130_fd_sc_hd__and2_4
  _1210_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[12] ),
    .X(_0761_)
  );


  sky130_fd_sc_hd__a21o_4
  _1211_
  (
    .A1(_0462_),
    .A2(\__uuf__._0027_ ),
    .B1(_0761_),
    .X(_0444_)
  );


  sky130_fd_sc_hd__and2_4
  _1212_
  (
    .A(shift),
    .B(\__uuf__._0029_ ),
    .X(_0762_)
  );


  sky130_fd_sc_hd__a21o_4
  _1213_
  (
    .A1(_0462_),
    .A2(\__uuf__._0025_ ),
    .B1(_0762_),
    .X(_0445_)
  );


  sky130_fd_sc_hd__and2_4
  _1214_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[11] ),
    .X(_0763_)
  );


  sky130_fd_sc_hd__a21o_4
  _1215_
  (
    .A1(_0462_),
    .A2(\__uuf__._0024_ ),
    .B1(_0763_),
    .X(_0446_)
  );


  sky130_fd_sc_hd__and2_4
  _1216_
  (
    .A(shift),
    .B(\__uuf__._0026_ ),
    .X(_0764_)
  );


  sky130_fd_sc_hd__a21o_4
  _1217_
  (
    .A1(_0462_),
    .A2(\__uuf__._0022_ ),
    .B1(_0764_),
    .X(_0447_)
  );


  sky130_fd_sc_hd__and2_4
  _1218_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[10] ),
    .X(_0765_)
  );


  sky130_fd_sc_hd__a21o_4
  _1219_
  (
    .A1(_0462_),
    .A2(\__uuf__._0021_ ),
    .B1(_0765_),
    .X(_0448_)
  );


  sky130_fd_sc_hd__and2_4
  _1220_
  (
    .A(shift),
    .B(\__uuf__._0023_ ),
    .X(_0766_)
  );


  sky130_fd_sc_hd__a21o_4
  _1221_
  (
    .A1(_0462_),
    .A2(\__uuf__._0019_ ),
    .B1(_0766_),
    .X(_0449_)
  );


  sky130_fd_sc_hd__and2_4
  _1222_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[9] ),
    .X(_0767_)
  );


  sky130_fd_sc_hd__a21o_4
  _1223_
  (
    .A1(_0462_),
    .A2(\__uuf__._0018_ ),
    .B1(_0767_),
    .X(_0450_)
  );


  sky130_fd_sc_hd__and2_4
  _1224_
  (
    .A(shift),
    .B(\__uuf__._0020_ ),
    .X(_0768_)
  );


  sky130_fd_sc_hd__a21o_4
  _1225_
  (
    .A1(_0462_),
    .A2(\__uuf__._0016_ ),
    .B1(_0768_),
    .X(_0451_)
  );


  sky130_fd_sc_hd__and2_4
  _1226_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[8] ),
    .X(_0769_)
  );


  sky130_fd_sc_hd__a21o_4
  _1227_
  (
    .A1(_0462_),
    .A2(\__uuf__._0015_ ),
    .B1(_0769_),
    .X(_0452_)
  );


  sky130_fd_sc_hd__and2_4
  _1228_
  (
    .A(shift),
    .B(\__uuf__._0017_ ),
    .X(_0770_)
  );


  sky130_fd_sc_hd__a21o_4
  _1229_
  (
    .A1(_0462_),
    .A2(\__uuf__._0013_ ),
    .B1(_0770_),
    .X(_0453_)
  );


  sky130_fd_sc_hd__and2_4
  _1230_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[7] ),
    .X(_0771_)
  );


  sky130_fd_sc_hd__a21o_4
  _1231_
  (
    .A1(_0462_),
    .A2(\__uuf__._0012_ ),
    .B1(_0771_),
    .X(_0454_)
  );


  sky130_fd_sc_hd__and2_4
  _1232_
  (
    .A(shift),
    .B(\__uuf__._0014_ ),
    .X(_0772_)
  );


  sky130_fd_sc_hd__a21o_4
  _1233_
  (
    .A1(_0462_),
    .A2(\__uuf__._0010_ ),
    .B1(_0772_),
    .X(_0455_)
  );


  sky130_fd_sc_hd__and2_4
  _1234_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[6] ),
    .X(_0773_)
  );


  sky130_fd_sc_hd__a21o_4
  _1235_
  (
    .A1(_0462_),
    .A2(\__uuf__._0009_ ),
    .B1(_0773_),
    .X(_0456_)
  );


  sky130_fd_sc_hd__and2_4
  _1236_
  (
    .A(shift),
    .B(\__uuf__._0011_ ),
    .X(_0774_)
  );


  sky130_fd_sc_hd__a21o_4
  _1237_
  (
    .A1(_0462_),
    .A2(\__uuf__._0007_ ),
    .B1(_0774_),
    .X(_0457_)
  );


  sky130_fd_sc_hd__and2_4
  _1238_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[5] ),
    .X(_0775_)
  );


  sky130_fd_sc_hd__a21o_4
  _1239_
  (
    .A1(_0462_),
    .A2(\__uuf__._0006_ ),
    .B1(_0775_),
    .X(_0458_)
  );


  sky130_fd_sc_hd__and2_4
  _1240_
  (
    .A(shift),
    .B(\__uuf__._0008_ ),
    .X(_0776_)
  );


  sky130_fd_sc_hd__a21o_4
  _1241_
  (
    .A1(_0462_),
    .A2(\__uuf__._0004_ ),
    .B1(_0776_),
    .X(_0459_)
  );


  sky130_fd_sc_hd__and2_4
  _1242_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[4] ),
    .X(_0777_)
  );


  sky130_fd_sc_hd__a21o_4
  _1243_
  (
    .A1(_0462_),
    .A2(\__uuf__._0003_ ),
    .B1(_0777_),
    .X(_0460_)
  );


  sky130_fd_sc_hd__and2_4
  _1244_
  (
    .A(shift),
    .B(\__uuf__._0005_ ),
    .X(_0778_)
  );


  sky130_fd_sc_hd__a21o_4
  _1245_
  (
    .A1(_0462_),
    .A2(\__uuf__._0001_ ),
    .B1(_0778_),
    .X(_0461_)
  );


  sky130_fd_sc_hd__and2_4
  _1246_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[3] ),
    .X(_0779_)
  );


  sky130_fd_sc_hd__a21o_4
  _1247_
  (
    .A1(_0462_),
    .A2(\__uuf__._0000_ ),
    .B1(_0779_),
    .X(_0260_)
  );


  sky130_fd_sc_hd__and2_4
  _1248_
  (
    .A(shift),
    .B(\__uuf__._0002_ ),
    .X(_0780_)
  );


  sky130_fd_sc_hd__a21o_4
  _1249_
  (
    .A1(_0462_),
    .A2(\__uuf__._0088_ ),
    .B1(_0780_),
    .X(_0261_)
  );


  sky130_fd_sc_hd__and2_4
  _1250_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[2] ),
    .X(_0781_)
  );


  sky130_fd_sc_hd__a21o_4
  _1251_
  (
    .A1(_0462_),
    .A2(\__uuf__._0087_ ),
    .B1(_0781_),
    .X(_0262_)
  );


  sky130_fd_sc_hd__and2_4
  _1252_
  (
    .A(shift),
    .B(\__uuf__._0089_ ),
    .X(_0782_)
  );


  sky130_fd_sc_hd__a21o_4
  _1253_
  (
    .A1(_0462_),
    .A2(\__uuf__._0085_ ),
    .B1(_0782_),
    .X(_0263_)
  );


  sky130_fd_sc_hd__and2_4
  _1254_
  (
    .A(shift),
    .B(\__uuf__.multiplier.csa0.y ),
    .X(_0783_)
  );


  sky130_fd_sc_hd__a21o_4
  _1255_
  (
    .A1(_0462_),
    .A2(\__uuf__._0084_ ),
    .B1(_0783_),
    .X(_0264_)
  );


  sky130_fd_sc_hd__and2_4
  _1256_
  (
    .A(shift),
    .B(\__uuf__._0086_ ),
    .X(_0784_)
  );


  sky130_fd_sc_hd__a21o_4
  _1257_
  (
    .A1(_0462_),
    .A2(\__uuf__._0092_ ),
    .B1(_0784_),
    .X(_0265_)
  );


  sky130_fd_sc_hd__and2_4
  _1258_
  (
    .A(shift),
    .B(\__uuf__.multiplier.pp[31] ),
    .X(_0785_)
  );


  sky130_fd_sc_hd__a21o_4
  _1259_
  (
    .A1(_0462_),
    .A2(\__uuf__._0093_ ),
    .B1(_0785_),
    .X(_0266_)
  );


  sky130_fd_sc_hd__and2_4
  _1260_
  (
    .A(shift),
    .B(\__uuf__.multiplier.tcmp.z ),
    .X(_0786_)
  );


  sky130_fd_sc_hd__a21o_4
  _1261_
  (
    .A1(_0462_),
    .A2(\__uuf__._0091_ ),
    .B1(_0786_),
    .X(_0267_)
  );


  sky130_fd_sc_hd__and2_4
  _1262_
  (
    .A(shift),
    .B(\__uuf__.multiplier.csa0.sum ),
    .X(_0787_)
  );


  sky130_fd_sc_hd__a21o_4
  _1263_
  (
    .A1(_0462_),
    .A2(\__uuf__._0090_ ),
    .B1(_0787_),
    .X(_0268_)
  );


  sky130_fd_sc_hd__and2_4
  _1264_
  (
    .A(shift),
    .B(\__uuf__.multiplier.csa0.sc ),
    .X(_0788_)
  );


  sky130_fd_sc_hd__a21o_4
  _1265_
  (
    .A1(_0462_),
    .A2(\__uuf__.fsm.newstate[0] ),
    .B1(_0788_),
    .X(_0269_)
  );


  sky130_fd_sc_hd__and2_4
  _1266_
  (
    .A(shift),
    .B(\__uuf__.fsm.state[0] ),
    .X(_0789_)
  );


  sky130_fd_sc_hd__a21o_4
  _1267_
  (
    .A1(_0462_),
    .A2(\__uuf__.fsm.newstate[1] ),
    .B1(_0789_),
    .X(_0270_)
  );


  sky130_fd_sc_hd__and2_4
  _1268_
  (
    .A(shift),
    .B(\__uuf__.fsm.state[1] ),
    .X(_0790_)
  );


  sky130_fd_sc_hd__a21o_4
  _1269_
  (
    .A1(_0462_),
    .A2(\__uuf__._0361_ ),
    .B1(_0790_),
    .X(_0271_)
  );


  sky130_fd_sc_hd__and2_4
  _1270_
  (
    .A(shift),
    .B(prod[0]),
    .X(_0791_)
  );


  sky130_fd_sc_hd__a21o_4
  _1271_
  (
    .A1(_0462_),
    .A2(\__uuf__._0362_ ),
    .B1(_0791_),
    .X(_0272_)
  );


  sky130_fd_sc_hd__and2_4
  _1272_
  (
    .A(shift),
    .B(prod[1]),
    .X(_0792_)
  );


  sky130_fd_sc_hd__a21o_4
  _1273_
  (
    .A1(_0462_),
    .A2(\__uuf__._0363_ ),
    .B1(_0792_),
    .X(_0273_)
  );


  sky130_fd_sc_hd__and2_4
  _1274_
  (
    .A(shift),
    .B(prod[2]),
    .X(_0793_)
  );


  sky130_fd_sc_hd__a21o_4
  _1275_
  (
    .A1(_0462_),
    .A2(\__uuf__._0364_ ),
    .B1(_0793_),
    .X(_0274_)
  );


  sky130_fd_sc_hd__and2_4
  _1276_
  (
    .A(shift),
    .B(prod[3]),
    .X(_0794_)
  );


  sky130_fd_sc_hd__a21o_4
  _1277_
  (
    .A1(_0462_),
    .A2(\__uuf__._0365_ ),
    .B1(_0794_),
    .X(_0275_)
  );


  sky130_fd_sc_hd__and2_4
  _1278_
  (
    .A(shift),
    .B(prod[4]),
    .X(_0795_)
  );


  sky130_fd_sc_hd__a21o_4
  _1279_
  (
    .A1(_0462_),
    .A2(\__uuf__._0366_ ),
    .B1(_0795_),
    .X(_0276_)
  );


  sky130_fd_sc_hd__and2_4
  _1280_
  (
    .A(shift),
    .B(prod[5]),
    .X(_0796_)
  );


  sky130_fd_sc_hd__a21o_4
  _1281_
  (
    .A1(_0462_),
    .A2(\__uuf__._0367_ ),
    .B1(_0796_),
    .X(_0277_)
  );


  sky130_fd_sc_hd__and2_4
  _1282_
  (
    .A(shift),
    .B(prod[6]),
    .X(_0797_)
  );


  sky130_fd_sc_hd__a21o_4
  _1283_
  (
    .A1(_0462_),
    .A2(\__uuf__._0368_ ),
    .B1(_0797_),
    .X(_0278_)
  );


  sky130_fd_sc_hd__and2_4
  _1284_
  (
    .A(shift),
    .B(prod[7]),
    .X(_0798_)
  );


  sky130_fd_sc_hd__a21o_4
  _1285_
  (
    .A1(_0462_),
    .A2(\__uuf__._0369_ ),
    .B1(_0798_),
    .X(_0279_)
  );


  sky130_fd_sc_hd__and2_4
  _1286_
  (
    .A(shift),
    .B(prod[8]),
    .X(_0799_)
  );


  sky130_fd_sc_hd__a21o_4
  _1287_
  (
    .A1(_0462_),
    .A2(\__uuf__._0370_ ),
    .B1(_0799_),
    .X(_0280_)
  );


  sky130_fd_sc_hd__and2_4
  _1288_
  (
    .A(shift),
    .B(prod[9]),
    .X(_0800_)
  );


  sky130_fd_sc_hd__a21o_4
  _1289_
  (
    .A1(_0462_),
    .A2(\__uuf__._0371_ ),
    .B1(_0800_),
    .X(_0281_)
  );


  sky130_fd_sc_hd__and2_4
  _1290_
  (
    .A(shift),
    .B(prod[10]),
    .X(_0801_)
  );


  sky130_fd_sc_hd__a21o_4
  _1291_
  (
    .A1(_0462_),
    .A2(\__uuf__._0372_ ),
    .B1(_0801_),
    .X(_0282_)
  );


  sky130_fd_sc_hd__and2_4
  _1292_
  (
    .A(shift),
    .B(prod[11]),
    .X(_0802_)
  );


  sky130_fd_sc_hd__a21o_4
  _1293_
  (
    .A1(_0462_),
    .A2(\__uuf__._0373_ ),
    .B1(_0802_),
    .X(_0283_)
  );


  sky130_fd_sc_hd__and2_4
  _1294_
  (
    .A(shift),
    .B(prod[12]),
    .X(_0803_)
  );


  sky130_fd_sc_hd__a21o_4
  _1295_
  (
    .A1(_0462_),
    .A2(\__uuf__._0374_ ),
    .B1(_0803_),
    .X(_0284_)
  );


  sky130_fd_sc_hd__and2_4
  _1296_
  (
    .A(shift),
    .B(prod[13]),
    .X(_0804_)
  );


  sky130_fd_sc_hd__a21o_4
  _1297_
  (
    .A1(_0462_),
    .A2(\__uuf__._0375_ ),
    .B1(_0804_),
    .X(_0285_)
  );


  sky130_fd_sc_hd__and2_4
  _1298_
  (
    .A(shift),
    .B(prod[14]),
    .X(_0805_)
  );


  sky130_fd_sc_hd__a21o_4
  _1299_
  (
    .A1(_0462_),
    .A2(\__uuf__._0376_ ),
    .B1(_0805_),
    .X(_0286_)
  );


  sky130_fd_sc_hd__and2_4
  _1300_
  (
    .A(shift),
    .B(prod[15]),
    .X(_0806_)
  );


  sky130_fd_sc_hd__a21o_4
  _1301_
  (
    .A1(_0462_),
    .A2(\__uuf__._0377_ ),
    .B1(_0806_),
    .X(_0287_)
  );


  sky130_fd_sc_hd__and2_4
  _1302_
  (
    .A(shift),
    .B(prod[16]),
    .X(_0807_)
  );


  sky130_fd_sc_hd__a21o_4
  _1303_
  (
    .A1(_0462_),
    .A2(\__uuf__._0378_ ),
    .B1(_0807_),
    .X(_0288_)
  );


  sky130_fd_sc_hd__and2_4
  _1304_
  (
    .A(shift),
    .B(prod[17]),
    .X(_0808_)
  );


  sky130_fd_sc_hd__a21o_4
  _1305_
  (
    .A1(_0462_),
    .A2(\__uuf__._0379_ ),
    .B1(_0808_),
    .X(_0289_)
  );


  sky130_fd_sc_hd__and2_4
  _1306_
  (
    .A(shift),
    .B(prod[18]),
    .X(_0809_)
  );


  sky130_fd_sc_hd__a21o_4
  _1307_
  (
    .A1(_0462_),
    .A2(\__uuf__._0380_ ),
    .B1(_0809_),
    .X(_0290_)
  );


  sky130_fd_sc_hd__and2_4
  _1308_
  (
    .A(shift),
    .B(prod[19]),
    .X(_0810_)
  );


  sky130_fd_sc_hd__a21o_4
  _1309_
  (
    .A1(_0462_),
    .A2(\__uuf__._0381_ ),
    .B1(_0810_),
    .X(_0291_)
  );


  sky130_fd_sc_hd__and2_4
  _1310_
  (
    .A(shift),
    .B(prod[20]),
    .X(_0811_)
  );


  sky130_fd_sc_hd__a21o_4
  _1311_
  (
    .A1(_0462_),
    .A2(\__uuf__._0382_ ),
    .B1(_0811_),
    .X(_0292_)
  );


  sky130_fd_sc_hd__and2_4
  _1312_
  (
    .A(shift),
    .B(prod[21]),
    .X(_0812_)
  );


  sky130_fd_sc_hd__a21o_4
  _1313_
  (
    .A1(_0462_),
    .A2(\__uuf__._0383_ ),
    .B1(_0812_),
    .X(_0293_)
  );


  sky130_fd_sc_hd__and2_4
  _1314_
  (
    .A(shift),
    .B(prod[22]),
    .X(_0813_)
  );


  sky130_fd_sc_hd__a21o_4
  _1315_
  (
    .A1(_0462_),
    .A2(\__uuf__._0384_ ),
    .B1(_0813_),
    .X(_0294_)
  );


  sky130_fd_sc_hd__and2_4
  _1316_
  (
    .A(shift),
    .B(prod[23]),
    .X(_0814_)
  );


  sky130_fd_sc_hd__a21o_4
  _1317_
  (
    .A1(_0462_),
    .A2(\__uuf__._0385_ ),
    .B1(_0814_),
    .X(_0295_)
  );


  sky130_fd_sc_hd__and2_4
  _1318_
  (
    .A(shift),
    .B(prod[24]),
    .X(_0815_)
  );


  sky130_fd_sc_hd__a21o_4
  _1319_
  (
    .A1(_0462_),
    .A2(\__uuf__._0386_ ),
    .B1(_0815_),
    .X(_0296_)
  );


  sky130_fd_sc_hd__and2_4
  _1320_
  (
    .A(shift),
    .B(prod[25]),
    .X(_0816_)
  );


  sky130_fd_sc_hd__a21o_4
  _1321_
  (
    .A1(_0462_),
    .A2(\__uuf__._0387_ ),
    .B1(_0816_),
    .X(_0297_)
  );


  sky130_fd_sc_hd__and2_4
  _1322_
  (
    .A(shift),
    .B(prod[26]),
    .X(_0817_)
  );


  sky130_fd_sc_hd__a21o_4
  _1323_
  (
    .A1(_0462_),
    .A2(\__uuf__._0388_ ),
    .B1(_0817_),
    .X(_0298_)
  );


  sky130_fd_sc_hd__and2_4
  _1324_
  (
    .A(shift),
    .B(prod[27]),
    .X(_0818_)
  );


  sky130_fd_sc_hd__a21o_4
  _1325_
  (
    .A1(_0462_),
    .A2(\__uuf__._0389_ ),
    .B1(_0818_),
    .X(_0299_)
  );


  sky130_fd_sc_hd__and2_4
  _1326_
  (
    .A(shift),
    .B(prod[28]),
    .X(_0819_)
  );


  sky130_fd_sc_hd__a21o_4
  _1327_
  (
    .A1(_0462_),
    .A2(\__uuf__._0390_ ),
    .B1(_0819_),
    .X(_0300_)
  );


  sky130_fd_sc_hd__and2_4
  _1328_
  (
    .A(shift),
    .B(prod[29]),
    .X(_0820_)
  );


  sky130_fd_sc_hd__a21o_4
  _1329_
  (
    .A1(_0462_),
    .A2(\__uuf__._0391_ ),
    .B1(_0820_),
    .X(_0301_)
  );


  sky130_fd_sc_hd__and2_4
  _1330_
  (
    .A(shift),
    .B(prod[30]),
    .X(_0821_)
  );


  sky130_fd_sc_hd__a21o_4
  _1331_
  (
    .A1(_0462_),
    .A2(\__uuf__._0392_ ),
    .B1(_0821_),
    .X(_0302_)
  );


  sky130_fd_sc_hd__and2_4
  _1332_
  (
    .A(shift),
    .B(prod[31]),
    .X(_0822_)
  );


  sky130_fd_sc_hd__a21o_4
  _1333_
  (
    .A1(_0462_),
    .A2(\__uuf__._0393_ ),
    .B1(_0822_),
    .X(_0303_)
  );


  sky130_fd_sc_hd__and2_4
  _1334_
  (
    .A(shift),
    .B(prod[32]),
    .X(_0823_)
  );


  sky130_fd_sc_hd__a21o_4
  _1335_
  (
    .A1(_0462_),
    .A2(\__uuf__._0394_ ),
    .B1(_0823_),
    .X(_0304_)
  );


  sky130_fd_sc_hd__and2_4
  _1336_
  (
    .A(shift),
    .B(prod[33]),
    .X(_0824_)
  );


  sky130_fd_sc_hd__a21o_4
  _1337_
  (
    .A1(_0462_),
    .A2(\__uuf__._0395_ ),
    .B1(_0824_),
    .X(_0305_)
  );


  sky130_fd_sc_hd__and2_4
  _1338_
  (
    .A(shift),
    .B(prod[34]),
    .X(_0825_)
  );


  sky130_fd_sc_hd__a21o_4
  _1339_
  (
    .A1(_0462_),
    .A2(\__uuf__._0396_ ),
    .B1(_0825_),
    .X(_0306_)
  );


  sky130_fd_sc_hd__and2_4
  _1340_
  (
    .A(shift),
    .B(prod[35]),
    .X(_0826_)
  );


  sky130_fd_sc_hd__a21o_4
  _1341_
  (
    .A1(_0462_),
    .A2(\__uuf__._0397_ ),
    .B1(_0826_),
    .X(_0307_)
  );


  sky130_fd_sc_hd__and2_4
  _1342_
  (
    .A(shift),
    .B(prod[36]),
    .X(_0827_)
  );


  sky130_fd_sc_hd__a21o_4
  _1343_
  (
    .A1(_0462_),
    .A2(\__uuf__._0398_ ),
    .B1(_0827_),
    .X(_0308_)
  );


  sky130_fd_sc_hd__and2_4
  _1344_
  (
    .A(shift),
    .B(prod[37]),
    .X(_0828_)
  );


  sky130_fd_sc_hd__a21o_4
  _1345_
  (
    .A1(_0462_),
    .A2(\__uuf__._0399_ ),
    .B1(_0828_),
    .X(_0309_)
  );


  sky130_fd_sc_hd__and2_4
  _1346_
  (
    .A(shift),
    .B(prod[38]),
    .X(_0829_)
  );


  sky130_fd_sc_hd__a21o_4
  _1347_
  (
    .A1(_0462_),
    .A2(\__uuf__._0400_ ),
    .B1(_0829_),
    .X(_0310_)
  );


  sky130_fd_sc_hd__and2_4
  _1348_
  (
    .A(shift),
    .B(prod[39]),
    .X(_0830_)
  );


  sky130_fd_sc_hd__a21o_4
  _1349_
  (
    .A1(_0462_),
    .A2(\__uuf__._0401_ ),
    .B1(_0830_),
    .X(_0311_)
  );


  sky130_fd_sc_hd__and2_4
  _1350_
  (
    .A(shift),
    .B(prod[40]),
    .X(_0831_)
  );


  sky130_fd_sc_hd__a21o_4
  _1351_
  (
    .A1(_0462_),
    .A2(\__uuf__._0402_ ),
    .B1(_0831_),
    .X(_0312_)
  );


  sky130_fd_sc_hd__and2_4
  _1352_
  (
    .A(shift),
    .B(prod[41]),
    .X(_0832_)
  );


  sky130_fd_sc_hd__a21o_4
  _1353_
  (
    .A1(_0462_),
    .A2(\__uuf__._0403_ ),
    .B1(_0832_),
    .X(_0313_)
  );


  sky130_fd_sc_hd__and2_4
  _1354_
  (
    .A(shift),
    .B(prod[42]),
    .X(_0833_)
  );


  sky130_fd_sc_hd__a21o_4
  _1355_
  (
    .A1(_0462_),
    .A2(\__uuf__._0404_ ),
    .B1(_0833_),
    .X(_0314_)
  );


  sky130_fd_sc_hd__and2_4
  _1356_
  (
    .A(shift),
    .B(prod[43]),
    .X(_0834_)
  );


  sky130_fd_sc_hd__a21o_4
  _1357_
  (
    .A1(_0462_),
    .A2(\__uuf__._0405_ ),
    .B1(_0834_),
    .X(_0315_)
  );


  sky130_fd_sc_hd__and2_4
  _1358_
  (
    .A(shift),
    .B(prod[44]),
    .X(_0835_)
  );


  sky130_fd_sc_hd__a21o_4
  _1359_
  (
    .A1(_0462_),
    .A2(\__uuf__._0406_ ),
    .B1(_0835_),
    .X(_0316_)
  );


  sky130_fd_sc_hd__and2_4
  _1360_
  (
    .A(shift),
    .B(prod[45]),
    .X(_0836_)
  );


  sky130_fd_sc_hd__a21o_4
  _1361_
  (
    .A1(_0462_),
    .A2(\__uuf__._0407_ ),
    .B1(_0836_),
    .X(_0317_)
  );


  sky130_fd_sc_hd__and2_4
  _1362_
  (
    .A(shift),
    .B(prod[46]),
    .X(_0837_)
  );


  sky130_fd_sc_hd__a21o_4
  _1363_
  (
    .A1(_0462_),
    .A2(\__uuf__._0408_ ),
    .B1(_0837_),
    .X(_0318_)
  );


  sky130_fd_sc_hd__and2_4
  _1364_
  (
    .A(shift),
    .B(prod[47]),
    .X(_0838_)
  );


  sky130_fd_sc_hd__a21o_4
  _1365_
  (
    .A1(_0462_),
    .A2(\__uuf__._0409_ ),
    .B1(_0838_),
    .X(_0319_)
  );


  sky130_fd_sc_hd__and2_4
  _1366_
  (
    .A(shift),
    .B(prod[48]),
    .X(_0839_)
  );


  sky130_fd_sc_hd__a21o_4
  _1367_
  (
    .A1(_0462_),
    .A2(\__uuf__._0410_ ),
    .B1(_0839_),
    .X(_0320_)
  );


  sky130_fd_sc_hd__and2_4
  _1368_
  (
    .A(shift),
    .B(prod[49]),
    .X(_0840_)
  );


  sky130_fd_sc_hd__a21o_4
  _1369_
  (
    .A1(_0462_),
    .A2(\__uuf__._0411_ ),
    .B1(_0840_),
    .X(_0321_)
  );


  sky130_fd_sc_hd__and2_4
  _1370_
  (
    .A(shift),
    .B(prod[50]),
    .X(_0841_)
  );


  sky130_fd_sc_hd__a21o_4
  _1371_
  (
    .A1(_0462_),
    .A2(\__uuf__._0412_ ),
    .B1(_0841_),
    .X(_0322_)
  );


  sky130_fd_sc_hd__and2_4
  _1372_
  (
    .A(shift),
    .B(prod[51]),
    .X(_0842_)
  );


  sky130_fd_sc_hd__a21o_4
  _1373_
  (
    .A1(_0462_),
    .A2(\__uuf__._0413_ ),
    .B1(_0842_),
    .X(_0323_)
  );


  sky130_fd_sc_hd__and2_4
  _1374_
  (
    .A(shift),
    .B(prod[52]),
    .X(_0843_)
  );


  sky130_fd_sc_hd__a21o_4
  _1375_
  (
    .A1(_0462_),
    .A2(\__uuf__._0414_ ),
    .B1(_0843_),
    .X(_0324_)
  );


  sky130_fd_sc_hd__and2_4
  _1376_
  (
    .A(shift),
    .B(prod[53]),
    .X(_0844_)
  );


  sky130_fd_sc_hd__a21o_4
  _1377_
  (
    .A1(_0462_),
    .A2(\__uuf__._0415_ ),
    .B1(_0844_),
    .X(_0325_)
  );


  sky130_fd_sc_hd__and2_4
  _1378_
  (
    .A(shift),
    .B(prod[54]),
    .X(_0845_)
  );


  sky130_fd_sc_hd__a21o_4
  _1379_
  (
    .A1(_0462_),
    .A2(\__uuf__._0416_ ),
    .B1(_0845_),
    .X(_0326_)
  );


  sky130_fd_sc_hd__and2_4
  _1380_
  (
    .A(shift),
    .B(prod[55]),
    .X(_0846_)
  );


  sky130_fd_sc_hd__a21o_4
  _1381_
  (
    .A1(_0462_),
    .A2(\__uuf__._0417_ ),
    .B1(_0846_),
    .X(_0327_)
  );


  sky130_fd_sc_hd__and2_4
  _1382_
  (
    .A(shift),
    .B(prod[56]),
    .X(_0847_)
  );


  sky130_fd_sc_hd__a21o_4
  _1383_
  (
    .A1(_0462_),
    .A2(\__uuf__._0418_ ),
    .B1(_0847_),
    .X(_0328_)
  );


  sky130_fd_sc_hd__and2_4
  _1384_
  (
    .A(shift),
    .B(prod[57]),
    .X(_0848_)
  );


  sky130_fd_sc_hd__a21o_4
  _1385_
  (
    .A1(_0462_),
    .A2(\__uuf__._0419_ ),
    .B1(_0848_),
    .X(_0329_)
  );


  sky130_fd_sc_hd__and2_4
  _1386_
  (
    .A(shift),
    .B(prod[58]),
    .X(_0849_)
  );


  sky130_fd_sc_hd__a21o_4
  _1387_
  (
    .A1(_0462_),
    .A2(\__uuf__._0420_ ),
    .B1(_0849_),
    .X(_0330_)
  );


  sky130_fd_sc_hd__and2_4
  _1388_
  (
    .A(shift),
    .B(prod[59]),
    .X(_0850_)
  );


  sky130_fd_sc_hd__a21o_4
  _1389_
  (
    .A1(_0462_),
    .A2(\__uuf__._0421_ ),
    .B1(_0850_),
    .X(_0331_)
  );


  sky130_fd_sc_hd__and2_4
  _1390_
  (
    .A(shift),
    .B(prod[60]),
    .X(_0851_)
  );


  sky130_fd_sc_hd__a21o_4
  _1391_
  (
    .A1(_0462_),
    .A2(\__uuf__._0422_ ),
    .B1(_0851_),
    .X(_0332_)
  );


  sky130_fd_sc_hd__and2_4
  _1392_
  (
    .A(shift),
    .B(prod[61]),
    .X(_0852_)
  );


  sky130_fd_sc_hd__a21o_4
  _1393_
  (
    .A1(_0462_),
    .A2(\__uuf__._0423_ ),
    .B1(_0852_),
    .X(_0333_)
  );


  sky130_fd_sc_hd__and2_4
  _1394_
  (
    .A(shift),
    .B(prod[62]),
    .X(_0853_)
  );


  sky130_fd_sc_hd__a21o_4
  _1395_
  (
    .A1(_0462_),
    .A2(\__uuf__._0424_ ),
    .B1(_0853_),
    .X(_0334_)
  );


  sky130_fd_sc_hd__and2_4
  _1396_
  (
    .A(shift),
    .B(prod[63]),
    .X(_0854_)
  );


  sky130_fd_sc_hd__a21o_4
  _1397_
  (
    .A1(_0462_),
    .A2(\__uuf__._0425_ ),
    .B1(_0854_),
    .X(_0335_)
  );


  sky130_fd_sc_hd__and2_4
  _1398_
  (
    .A(shift),
    .B(\__uuf__.count[0] ),
    .X(_0855_)
  );


  sky130_fd_sc_hd__a21o_4
  _1399_
  (
    .A1(_0462_),
    .A2(\__uuf__._0426_ ),
    .B1(_0855_),
    .X(_0336_)
  );


  sky130_fd_sc_hd__and2_4
  _1400_
  (
    .A(shift),
    .B(\__uuf__.count[1] ),
    .X(_0856_)
  );


  sky130_fd_sc_hd__a21o_4
  _1401_
  (
    .A1(_0462_),
    .A2(\__uuf__._0427_ ),
    .B1(_0856_),
    .X(_0337_)
  );


  sky130_fd_sc_hd__and2_4
  _1402_
  (
    .A(shift),
    .B(\__uuf__.count[2] ),
    .X(_0857_)
  );


  sky130_fd_sc_hd__a21o_4
  _1403_
  (
    .A1(_0462_),
    .A2(\__uuf__._0428_ ),
    .B1(_0857_),
    .X(_0338_)
  );


  sky130_fd_sc_hd__and2_4
  _1404_
  (
    .A(shift),
    .B(\__uuf__.count[3] ),
    .X(_0858_)
  );


  sky130_fd_sc_hd__a21o_4
  _1405_
  (
    .A1(_0462_),
    .A2(\__uuf__._0429_ ),
    .B1(_0858_),
    .X(_0339_)
  );


  sky130_fd_sc_hd__and2_4
  _1406_
  (
    .A(shift),
    .B(\__uuf__.count[4] ),
    .X(_0859_)
  );


  sky130_fd_sc_hd__a21o_4
  _1407_
  (
    .A1(_0462_),
    .A2(\__uuf__._0430_ ),
    .B1(_0859_),
    .X(_0340_)
  );


  sky130_fd_sc_hd__and2_4
  _1408_
  (
    .A(shift),
    .B(\__uuf__.count[5] ),
    .X(_0860_)
  );


  sky130_fd_sc_hd__a21o_4
  _1409_
  (
    .A1(_0462_),
    .A2(\__uuf__._0431_ ),
    .B1(_0860_),
    .X(_0341_)
  );


  sky130_fd_sc_hd__and2_4
  _1410_
  (
    .A(test),
    .B(tck),
    .X(_0861_)
  );


  sky130_fd_sc_hd__a21o_4
  _1411_
  (
    .A1(_0463_),
    .A2(clk),
    .B1(_0861_),
    .X(\__uuf__.__clk_source__ )
  );


  sky130_fd_sc_hd__inv_2
  _1412_
  (
    .A(rst),
    .Y(_0127_)
  );


  sky130_fd_sc_hd__inv_2
  _1413_
  (
    .A(rst),
    .Y(_0126_)
  );


  sky130_fd_sc_hd__inv_2
  _1414_
  (
    .A(rst),
    .Y(_0125_)
  );


  sky130_fd_sc_hd__inv_2
  _1415_
  (
    .A(rst),
    .Y(_0124_)
  );


  sky130_fd_sc_hd__inv_2
  _1416_
  (
    .A(rst),
    .Y(_0123_)
  );


  sky130_fd_sc_hd__inv_2
  _1417_
  (
    .A(rst),
    .Y(_0122_)
  );


  sky130_fd_sc_hd__inv_2
  _1418_
  (
    .A(rst),
    .Y(_0121_)
  );


  sky130_fd_sc_hd__inv_2
  _1419_
  (
    .A(rst),
    .Y(_0120_)
  );


  sky130_fd_sc_hd__inv_2
  _1420_
  (
    .A(rst),
    .Y(_0119_)
  );


  sky130_fd_sc_hd__inv_2
  _1421_
  (
    .A(rst),
    .Y(_0118_)
  );


  sky130_fd_sc_hd__inv_2
  _1422_
  (
    .A(rst),
    .Y(_0117_)
  );


  sky130_fd_sc_hd__inv_2
  _1423_
  (
    .A(rst),
    .Y(_0116_)
  );


  sky130_fd_sc_hd__inv_2
  _1424_
  (
    .A(rst),
    .Y(_0115_)
  );


  sky130_fd_sc_hd__inv_2
  _1425_
  (
    .A(rst),
    .Y(_0114_)
  );


  sky130_fd_sc_hd__inv_2
  _1426_
  (
    .A(rst),
    .Y(_0113_)
  );


  sky130_fd_sc_hd__inv_2
  _1427_
  (
    .A(rst),
    .Y(_0112_)
  );


  sky130_fd_sc_hd__inv_2
  _1428_
  (
    .A(rst),
    .Y(_0111_)
  );


  sky130_fd_sc_hd__inv_2
  _1429_
  (
    .A(rst),
    .Y(_0110_)
  );


  sky130_fd_sc_hd__inv_2
  _1430_
  (
    .A(rst),
    .Y(_0109_)
  );


  sky130_fd_sc_hd__inv_2
  _1431_
  (
    .A(rst),
    .Y(_0108_)
  );


  sky130_fd_sc_hd__inv_2
  _1432_
  (
    .A(rst),
    .Y(_0107_)
  );


  sky130_fd_sc_hd__inv_2
  _1433_
  (
    .A(rst),
    .Y(_0106_)
  );


  sky130_fd_sc_hd__inv_2
  _1434_
  (
    .A(rst),
    .Y(_0105_)
  );


  sky130_fd_sc_hd__inv_2
  _1435_
  (
    .A(rst),
    .Y(_0104_)
  );


  sky130_fd_sc_hd__inv_2
  _1436_
  (
    .A(rst),
    .Y(_0103_)
  );


  sky130_fd_sc_hd__inv_2
  _1437_
  (
    .A(rst),
    .Y(_0102_)
  );


  sky130_fd_sc_hd__inv_2
  _1438_
  (
    .A(rst),
    .Y(_0101_)
  );


  sky130_fd_sc_hd__inv_2
  _1439_
  (
    .A(rst),
    .Y(_0100_)
  );


  sky130_fd_sc_hd__inv_2
  _1440_
  (
    .A(rst),
    .Y(_0099_)
  );


  sky130_fd_sc_hd__inv_2
  _1441_
  (
    .A(rst),
    .Y(_0098_)
  );


  sky130_fd_sc_hd__inv_2
  _1442_
  (
    .A(rst),
    .Y(_0097_)
  );


  sky130_fd_sc_hd__inv_2
  _1443_
  (
    .A(rst),
    .Y(_0096_)
  );


  sky130_fd_sc_hd__inv_2
  _1444_
  (
    .A(rst),
    .Y(_0095_)
  );


  sky130_fd_sc_hd__inv_2
  _1445_
  (
    .A(rst),
    .Y(_0094_)
  );


  sky130_fd_sc_hd__inv_2
  _1446_
  (
    .A(rst),
    .Y(_0093_)
  );


  sky130_fd_sc_hd__inv_2
  _1447_
  (
    .A(rst),
    .Y(_0092_)
  );


  sky130_fd_sc_hd__inv_2
  _1448_
  (
    .A(rst),
    .Y(_0091_)
  );


  sky130_fd_sc_hd__inv_2
  _1449_
  (
    .A(rst),
    .Y(_0090_)
  );


  sky130_fd_sc_hd__inv_2
  _1450_
  (
    .A(rst),
    .Y(_0089_)
  );


  sky130_fd_sc_hd__inv_2
  _1451_
  (
    .A(rst),
    .Y(_0088_)
  );


  sky130_fd_sc_hd__inv_2
  _1452_
  (
    .A(rst),
    .Y(_0087_)
  );


  sky130_fd_sc_hd__inv_2
  _1453_
  (
    .A(rst),
    .Y(_0086_)
  );


  sky130_fd_sc_hd__inv_2
  _1454_
  (
    .A(rst),
    .Y(_0085_)
  );


  sky130_fd_sc_hd__inv_2
  _1455_
  (
    .A(rst),
    .Y(_0084_)
  );


  sky130_fd_sc_hd__inv_2
  _1456_
  (
    .A(rst),
    .Y(_0083_)
  );


  sky130_fd_sc_hd__inv_2
  _1457_
  (
    .A(rst),
    .Y(_0082_)
  );


  sky130_fd_sc_hd__inv_2
  _1458_
  (
    .A(rst),
    .Y(_0081_)
  );


  sky130_fd_sc_hd__inv_2
  _1459_
  (
    .A(rst),
    .Y(_0080_)
  );


  sky130_fd_sc_hd__inv_2
  _1460_
  (
    .A(rst),
    .Y(_0079_)
  );


  sky130_fd_sc_hd__inv_2
  _1461_
  (
    .A(rst),
    .Y(_0078_)
  );


  sky130_fd_sc_hd__inv_2
  _1462_
  (
    .A(rst),
    .Y(_0077_)
  );


  sky130_fd_sc_hd__inv_2
  _1463_
  (
    .A(rst),
    .Y(_0076_)
  );


  sky130_fd_sc_hd__inv_2
  _1464_
  (
    .A(rst),
    .Y(_0075_)
  );


  sky130_fd_sc_hd__inv_2
  _1465_
  (
    .A(rst),
    .Y(_0074_)
  );


  sky130_fd_sc_hd__inv_2
  _1466_
  (
    .A(rst),
    .Y(_0073_)
  );


  sky130_fd_sc_hd__inv_2
  _1467_
  (
    .A(rst),
    .Y(_0072_)
  );


  sky130_fd_sc_hd__inv_2
  _1468_
  (
    .A(rst),
    .Y(_0071_)
  );


  sky130_fd_sc_hd__inv_2
  _1469_
  (
    .A(rst),
    .Y(_0070_)
  );


  sky130_fd_sc_hd__inv_2
  _1470_
  (
    .A(rst),
    .Y(_0069_)
  );


  sky130_fd_sc_hd__inv_2
  _1471_
  (
    .A(rst),
    .Y(_0068_)
  );


  sky130_fd_sc_hd__inv_2
  _1472_
  (
    .A(rst),
    .Y(_0067_)
  );


  sky130_fd_sc_hd__inv_2
  _1473_
  (
    .A(rst),
    .Y(_0066_)
  );


  sky130_fd_sc_hd__inv_2
  _1474_
  (
    .A(rst),
    .Y(_0065_)
  );


  sky130_fd_sc_hd__inv_2
  _1475_
  (
    .A(rst),
    .Y(_0064_)
  );


  sky130_fd_sc_hd__inv_2
  _1476_
  (
    .A(rst),
    .Y(_0063_)
  );


  sky130_fd_sc_hd__inv_2
  _1477_
  (
    .A(rst),
    .Y(_0062_)
  );


  sky130_fd_sc_hd__inv_2
  _1478_
  (
    .A(rst),
    .Y(_0061_)
  );


  sky130_fd_sc_hd__inv_2
  _1479_
  (
    .A(rst),
    .Y(_0060_)
  );


  sky130_fd_sc_hd__inv_2
  _1480_
  (
    .A(rst),
    .Y(_0059_)
  );


  sky130_fd_sc_hd__inv_2
  _1481_
  (
    .A(rst),
    .Y(_0058_)
  );


  sky130_fd_sc_hd__inv_2
  _1482_
  (
    .A(rst),
    .Y(_0057_)
  );


  sky130_fd_sc_hd__inv_2
  _1483_
  (
    .A(rst),
    .Y(_0056_)
  );


  sky130_fd_sc_hd__inv_2
  _1484_
  (
    .A(rst),
    .Y(_0055_)
  );


  sky130_fd_sc_hd__inv_2
  _1485_
  (
    .A(rst),
    .Y(_0054_)
  );


  sky130_fd_sc_hd__inv_2
  _1486_
  (
    .A(rst),
    .Y(_0053_)
  );


  sky130_fd_sc_hd__inv_2
  _1487_
  (
    .A(rst),
    .Y(_0052_)
  );


  sky130_fd_sc_hd__inv_2
  _1488_
  (
    .A(rst),
    .Y(_0051_)
  );


  sky130_fd_sc_hd__inv_2
  _1489_
  (
    .A(rst),
    .Y(_0050_)
  );


  sky130_fd_sc_hd__inv_2
  _1490_
  (
    .A(rst),
    .Y(_0049_)
  );


  sky130_fd_sc_hd__inv_2
  _1491_
  (
    .A(rst),
    .Y(_0048_)
  );


  sky130_fd_sc_hd__inv_2
  _1492_
  (
    .A(rst),
    .Y(_0047_)
  );


  sky130_fd_sc_hd__inv_2
  _1493_
  (
    .A(rst),
    .Y(_0046_)
  );


  sky130_fd_sc_hd__inv_2
  _1494_
  (
    .A(rst),
    .Y(_0045_)
  );


  sky130_fd_sc_hd__inv_2
  _1495_
  (
    .A(rst),
    .Y(_0044_)
  );


  sky130_fd_sc_hd__inv_2
  _1496_
  (
    .A(rst),
    .Y(_0043_)
  );


  sky130_fd_sc_hd__inv_2
  _1497_
  (
    .A(rst),
    .Y(_0042_)
  );


  sky130_fd_sc_hd__inv_2
  _1498_
  (
    .A(rst),
    .Y(_0041_)
  );


  sky130_fd_sc_hd__inv_2
  _1499_
  (
    .A(rst),
    .Y(_0040_)
  );


  sky130_fd_sc_hd__inv_2
  _1500_
  (
    .A(rst),
    .Y(_0039_)
  );


  sky130_fd_sc_hd__inv_2
  _1501_
  (
    .A(rst),
    .Y(_0038_)
  );


  sky130_fd_sc_hd__inv_2
  _1502_
  (
    .A(rst),
    .Y(_0037_)
  );


  sky130_fd_sc_hd__inv_2
  _1503_
  (
    .A(rst),
    .Y(_0036_)
  );


  sky130_fd_sc_hd__inv_2
  _1504_
  (
    .A(rst),
    .Y(_0035_)
  );


  sky130_fd_sc_hd__inv_2
  _1505_
  (
    .A(rst),
    .Y(_0034_)
  );


  sky130_fd_sc_hd__inv_2
  _1506_
  (
    .A(rst),
    .Y(_0033_)
  );


  sky130_fd_sc_hd__inv_2
  _1507_
  (
    .A(rst),
    .Y(_0032_)
  );


  sky130_fd_sc_hd__inv_2
  _1508_
  (
    .A(rst),
    .Y(_0031_)
  );


  sky130_fd_sc_hd__inv_2
  _1509_
  (
    .A(rst),
    .Y(_0030_)
  );


  sky130_fd_sc_hd__inv_2
  _1510_
  (
    .A(rst),
    .Y(_0029_)
  );


  sky130_fd_sc_hd__inv_2
  _1511_
  (
    .A(rst),
    .Y(_0028_)
  );


  sky130_fd_sc_hd__inv_2
  _1512_
  (
    .A(rst),
    .Y(_0027_)
  );


  sky130_fd_sc_hd__inv_2
  _1513_
  (
    .A(rst),
    .Y(_0026_)
  );


  sky130_fd_sc_hd__inv_2
  _1514_
  (
    .A(rst),
    .Y(_0025_)
  );


  sky130_fd_sc_hd__inv_2
  _1515_
  (
    .A(rst),
    .Y(_0024_)
  );


  sky130_fd_sc_hd__inv_2
  _1516_
  (
    .A(rst),
    .Y(_0023_)
  );


  sky130_fd_sc_hd__inv_2
  _1517_
  (
    .A(rst),
    .Y(_0022_)
  );


  sky130_fd_sc_hd__inv_2
  _1518_
  (
    .A(rst),
    .Y(_0021_)
  );


  sky130_fd_sc_hd__inv_2
  _1519_
  (
    .A(rst),
    .Y(_0020_)
  );


  sky130_fd_sc_hd__inv_2
  _1520_
  (
    .A(rst),
    .Y(_0019_)
  );


  sky130_fd_sc_hd__inv_2
  _1521_
  (
    .A(rst),
    .Y(_0018_)
  );


  sky130_fd_sc_hd__inv_2
  _1522_
  (
    .A(rst),
    .Y(_0017_)
  );


  sky130_fd_sc_hd__inv_2
  _1523_
  (
    .A(rst),
    .Y(_0016_)
  );


  sky130_fd_sc_hd__inv_2
  _1524_
  (
    .A(rst),
    .Y(_0015_)
  );


  sky130_fd_sc_hd__inv_2
  _1525_
  (
    .A(rst),
    .Y(_0014_)
  );


  sky130_fd_sc_hd__inv_2
  _1526_
  (
    .A(rst),
    .Y(_0013_)
  );


  sky130_fd_sc_hd__inv_2
  _1527_
  (
    .A(rst),
    .Y(_0012_)
  );


  sky130_fd_sc_hd__inv_2
  _1528_
  (
    .A(rst),
    .Y(_0011_)
  );


  sky130_fd_sc_hd__inv_2
  _1529_
  (
    .A(rst),
    .Y(_0010_)
  );


  sky130_fd_sc_hd__inv_2
  _1530_
  (
    .A(rst),
    .Y(_0009_)
  );


  sky130_fd_sc_hd__inv_2
  _1531_
  (
    .A(rst),
    .Y(_0008_)
  );


  sky130_fd_sc_hd__inv_2
  _1532_
  (
    .A(rst),
    .Y(_0007_)
  );


  sky130_fd_sc_hd__inv_2
  _1533_
  (
    .A(rst),
    .Y(_0006_)
  );


  sky130_fd_sc_hd__inv_2
  _1534_
  (
    .A(rst),
    .Y(_0005_)
  );


  sky130_fd_sc_hd__inv_2
  _1535_
  (
    .A(rst),
    .Y(_0004_)
  );


  sky130_fd_sc_hd__inv_2
  _1536_
  (
    .A(rst),
    .Y(_0003_)
  );


  sky130_fd_sc_hd__inv_2
  _1537_
  (
    .A(rst),
    .Y(_0002_)
  );


  sky130_fd_sc_hd__inv_2
  _1538_
  (
    .A(rst),
    .Y(_0001_)
  );


  sky130_fd_sc_hd__inv_2
  _1539_
  (
    .A(rst),
    .Y(_0000_)
  );


  sky130_fd_sc_hd__inv_2
  _1540_
  (
    .A(rst),
    .Y(_0129_)
  );


  sky130_fd_sc_hd__inv_2
  _1541_
  (
    .A(rst),
    .Y(_0128_)
  );


  sky130_fd_sc_hd__inv_2
  _1542_
  (
    .A(shift),
    .Y(_0462_)
  );


  sky130_fd_sc_hd__inv_2
  _1543_
  (
    .A(test),
    .Y(_0463_)
  );


  sky130_fd_sc_hd__and2_4
  _1544_
  (
    .A(\__BoundaryScanRegister_input_0__.sout ),
    .B(test),
    .X(_0464_)
  );


  sky130_fd_sc_hd__a21o_4
  _1545_
  (
    .A1(mc[0]),
    .A2(_0463_),
    .B1(_0464_),
    .X(\__BoundaryScanRegister_input_0__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1546_
  (
    .A(sin),
    .B(shift),
    .X(_0465_)
  );


  sky130_fd_sc_hd__a21o_4
  _1547_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_0__.dout ),
    .B1(_0465_),
    .X(_0130_)
  );


  sky130_fd_sc_hd__and2_4
  _1548_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_10__.sout ),
    .X(_0466_)
  );


  sky130_fd_sc_hd__a21o_4
  _1549_
  (
    .A1(_0463_),
    .A2(mc[10]),
    .B1(_0466_),
    .X(\__BoundaryScanRegister_input_10__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1550_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_10__.sin ),
    .X(_0467_)
  );


  sky130_fd_sc_hd__a21o_4
  _1551_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_10__.dout ),
    .B1(_0467_),
    .X(_0131_)
  );


  sky130_fd_sc_hd__and2_4
  _1552_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_11__.sout ),
    .X(_0468_)
  );


  sky130_fd_sc_hd__a21o_4
  _1553_
  (
    .A1(_0463_),
    .A2(mc[11]),
    .B1(_0468_),
    .X(\__BoundaryScanRegister_input_11__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1554_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_10__.sout ),
    .X(_0469_)
  );


  sky130_fd_sc_hd__a21o_4
  _1555_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_11__.dout ),
    .B1(_0469_),
    .X(_0132_)
  );


  sky130_fd_sc_hd__and2_4
  _1556_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_12__.sout ),
    .X(_0470_)
  );


  sky130_fd_sc_hd__a21o_4
  _1557_
  (
    .A1(_0463_),
    .A2(mc[12]),
    .B1(_0470_),
    .X(\__BoundaryScanRegister_input_12__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1558_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_11__.sout ),
    .X(_0471_)
  );


  sky130_fd_sc_hd__a21o_4
  _1559_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_12__.dout ),
    .B1(_0471_),
    .X(_0133_)
  );


  sky130_fd_sc_hd__and2_4
  _1560_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_13__.sout ),
    .X(_0472_)
  );


  sky130_fd_sc_hd__a21o_4
  _1561_
  (
    .A1(_0463_),
    .A2(mc[13]),
    .B1(_0472_),
    .X(\__BoundaryScanRegister_input_13__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1562_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_12__.sout ),
    .X(_0473_)
  );


  sky130_fd_sc_hd__a21o_4
  _1563_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_13__.dout ),
    .B1(_0473_),
    .X(_0134_)
  );


  sky130_fd_sc_hd__and2_4
  _1564_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_14__.sout ),
    .X(_0474_)
  );


  sky130_fd_sc_hd__a21o_4
  _1565_
  (
    .A1(_0463_),
    .A2(mc[14]),
    .B1(_0474_),
    .X(\__BoundaryScanRegister_input_14__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1566_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_13__.sout ),
    .X(_0475_)
  );


  sky130_fd_sc_hd__a21o_4
  _1567_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_14__.dout ),
    .B1(_0475_),
    .X(_0135_)
  );


  sky130_fd_sc_hd__and2_4
  _1568_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_15__.sout ),
    .X(_0476_)
  );


  sky130_fd_sc_hd__a21o_4
  _1569_
  (
    .A1(_0463_),
    .A2(mc[15]),
    .B1(_0476_),
    .X(\__BoundaryScanRegister_input_15__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1570_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_14__.sout ),
    .X(_0477_)
  );


  sky130_fd_sc_hd__a21o_4
  _1571_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_15__.dout ),
    .B1(_0477_),
    .X(_0136_)
  );


  sky130_fd_sc_hd__and2_4
  _1572_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_16__.sout ),
    .X(_0478_)
  );


  sky130_fd_sc_hd__a21o_4
  _1573_
  (
    .A1(_0463_),
    .A2(mc[16]),
    .B1(_0478_),
    .X(\__BoundaryScanRegister_input_16__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1574_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_15__.sout ),
    .X(_0479_)
  );


  sky130_fd_sc_hd__a21o_4
  _1575_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_16__.dout ),
    .B1(_0479_),
    .X(_0137_)
  );


  sky130_fd_sc_hd__and2_4
  _1576_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_17__.sout ),
    .X(_0480_)
  );


  sky130_fd_sc_hd__a21o_4
  _1577_
  (
    .A1(_0463_),
    .A2(mc[17]),
    .B1(_0480_),
    .X(\__BoundaryScanRegister_input_17__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1578_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_16__.sout ),
    .X(_0481_)
  );


  sky130_fd_sc_hd__a21o_4
  _1579_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_17__.dout ),
    .B1(_0481_),
    .X(_0138_)
  );


  sky130_fd_sc_hd__and2_4
  _1580_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_18__.sout ),
    .X(_0482_)
  );


  sky130_fd_sc_hd__a21o_4
  _1581_
  (
    .A1(_0463_),
    .A2(mc[18]),
    .B1(_0482_),
    .X(\__BoundaryScanRegister_input_18__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1582_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_17__.sout ),
    .X(_0483_)
  );


  sky130_fd_sc_hd__a21o_4
  _1583_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_18__.dout ),
    .B1(_0483_),
    .X(_0139_)
  );


  sky130_fd_sc_hd__and2_4
  _1584_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_19__.sout ),
    .X(_0484_)
  );


  sky130_fd_sc_hd__a21o_4
  _1585_
  (
    .A1(_0463_),
    .A2(mc[19]),
    .B1(_0484_),
    .X(\__BoundaryScanRegister_input_19__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1586_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_18__.sout ),
    .X(_0485_)
  );


  sky130_fd_sc_hd__a21o_4
  _1587_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_19__.dout ),
    .B1(_0485_),
    .X(_0140_)
  );


  sky130_fd_sc_hd__and2_4
  _1588_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_1__.sout ),
    .X(_0486_)
  );


  sky130_fd_sc_hd__a21o_4
  _1589_
  (
    .A1(_0463_),
    .A2(mc[1]),
    .B1(_0486_),
    .X(\__BoundaryScanRegister_input_1__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1590_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_0__.sout ),
    .X(_0487_)
  );


  sky130_fd_sc_hd__a21o_4
  _1591_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_1__.dout ),
    .B1(_0487_),
    .X(_0141_)
  );


  sky130_fd_sc_hd__and2_4
  _1592_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_20__.sout ),
    .X(_0488_)
  );


  sky130_fd_sc_hd__a21o_4
  _1593_
  (
    .A1(_0463_),
    .A2(mc[20]),
    .B1(_0488_),
    .X(\__BoundaryScanRegister_input_20__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1594_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_19__.sout ),
    .X(_0489_)
  );


  sky130_fd_sc_hd__a21o_4
  _1595_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_20__.dout ),
    .B1(_0489_),
    .X(_0142_)
  );


  sky130_fd_sc_hd__and2_4
  _1596_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_21__.sout ),
    .X(_0490_)
  );


  sky130_fd_sc_hd__a21o_4
  _1597_
  (
    .A1(_0463_),
    .A2(mc[21]),
    .B1(_0490_),
    .X(\__BoundaryScanRegister_input_21__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1598_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_20__.sout ),
    .X(_0491_)
  );


  sky130_fd_sc_hd__a21o_4
  _1599_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_21__.dout ),
    .B1(_0491_),
    .X(_0143_)
  );


  sky130_fd_sc_hd__and2_4
  _1600_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_22__.sout ),
    .X(_0492_)
  );


  sky130_fd_sc_hd__a21o_4
  _1601_
  (
    .A1(_0463_),
    .A2(mc[22]),
    .B1(_0492_),
    .X(\__BoundaryScanRegister_input_22__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1602_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_21__.sout ),
    .X(_0493_)
  );


  sky130_fd_sc_hd__a21o_4
  _1603_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_22__.dout ),
    .B1(_0493_),
    .X(_0144_)
  );


  sky130_fd_sc_hd__and2_4
  _1604_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_23__.sout ),
    .X(_0494_)
  );


  sky130_fd_sc_hd__a21o_4
  _1605_
  (
    .A1(_0463_),
    .A2(mc[23]),
    .B1(_0494_),
    .X(\__BoundaryScanRegister_input_23__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1606_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_22__.sout ),
    .X(_0495_)
  );


  sky130_fd_sc_hd__a21o_4
  _1607_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_23__.dout ),
    .B1(_0495_),
    .X(_0145_)
  );


  sky130_fd_sc_hd__and2_4
  _1608_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_24__.sout ),
    .X(_0496_)
  );


  sky130_fd_sc_hd__a21o_4
  _1609_
  (
    .A1(_0463_),
    .A2(mc[24]),
    .B1(_0496_),
    .X(\__BoundaryScanRegister_input_24__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1610_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_23__.sout ),
    .X(_0497_)
  );


  sky130_fd_sc_hd__a21o_4
  _1611_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_24__.dout ),
    .B1(_0497_),
    .X(_0146_)
  );


  sky130_fd_sc_hd__and2_4
  _1612_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_25__.sout ),
    .X(_0498_)
  );


  sky130_fd_sc_hd__a21o_4
  _1613_
  (
    .A1(_0463_),
    .A2(mc[25]),
    .B1(_0498_),
    .X(\__BoundaryScanRegister_input_25__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1614_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_24__.sout ),
    .X(_0499_)
  );


  sky130_fd_sc_hd__a21o_4
  _1615_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_25__.dout ),
    .B1(_0499_),
    .X(_0147_)
  );


  sky130_fd_sc_hd__and2_4
  _1616_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_26__.sout ),
    .X(_0500_)
  );


  sky130_fd_sc_hd__a21o_4
  _1617_
  (
    .A1(_0463_),
    .A2(mc[26]),
    .B1(_0500_),
    .X(\__BoundaryScanRegister_input_26__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1618_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_25__.sout ),
    .X(_0501_)
  );


  sky130_fd_sc_hd__a21o_4
  _1619_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_26__.dout ),
    .B1(_0501_),
    .X(_0148_)
  );


  sky130_fd_sc_hd__and2_4
  _1620_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_27__.sout ),
    .X(_0502_)
  );


  sky130_fd_sc_hd__a21o_4
  _1621_
  (
    .A1(_0463_),
    .A2(mc[27]),
    .B1(_0502_),
    .X(\__BoundaryScanRegister_input_27__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1622_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_26__.sout ),
    .X(_0503_)
  );


  sky130_fd_sc_hd__a21o_4
  _1623_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_27__.dout ),
    .B1(_0503_),
    .X(_0149_)
  );


  sky130_fd_sc_hd__and2_4
  _1624_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_28__.sout ),
    .X(_0504_)
  );


  sky130_fd_sc_hd__a21o_4
  _1625_
  (
    .A1(_0463_),
    .A2(mc[28]),
    .B1(_0504_),
    .X(\__BoundaryScanRegister_input_28__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1626_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_27__.sout ),
    .X(_0505_)
  );


  sky130_fd_sc_hd__a21o_4
  _1627_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_28__.dout ),
    .B1(_0505_),
    .X(_0150_)
  );


  sky130_fd_sc_hd__and2_4
  _1628_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_29__.sout ),
    .X(_0506_)
  );


  sky130_fd_sc_hd__a21o_4
  _1629_
  (
    .A1(_0463_),
    .A2(mc[29]),
    .B1(_0506_),
    .X(\__BoundaryScanRegister_input_29__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1630_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_28__.sout ),
    .X(_0507_)
  );


  sky130_fd_sc_hd__a21o_4
  _1631_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_29__.dout ),
    .B1(_0507_),
    .X(_0151_)
  );


  sky130_fd_sc_hd__and2_4
  _1632_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_2__.sout ),
    .X(_0508_)
  );


  sky130_fd_sc_hd__a21o_4
  _1633_
  (
    .A1(_0463_),
    .A2(mc[2]),
    .B1(_0508_),
    .X(\__BoundaryScanRegister_input_2__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1634_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_1__.sout ),
    .X(_0509_)
  );


  sky130_fd_sc_hd__a21o_4
  _1635_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_2__.dout ),
    .B1(_0509_),
    .X(_0152_)
  );


  sky130_fd_sc_hd__and2_4
  _1636_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_30__.sout ),
    .X(_0510_)
  );


  sky130_fd_sc_hd__a21o_4
  _1637_
  (
    .A1(_0463_),
    .A2(mc[30]),
    .B1(_0510_),
    .X(\__BoundaryScanRegister_input_30__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1638_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_29__.sout ),
    .X(_0511_)
  );


  sky130_fd_sc_hd__a21o_4
  _1639_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_30__.dout ),
    .B1(_0511_),
    .X(_0153_)
  );


  sky130_fd_sc_hd__and2_4
  _1640_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_31__.sout ),
    .X(_0512_)
  );


  sky130_fd_sc_hd__a21o_4
  _1641_
  (
    .A1(_0463_),
    .A2(mc[31]),
    .B1(_0512_),
    .X(\__BoundaryScanRegister_input_31__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1642_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_30__.sout ),
    .X(_0513_)
  );


  sky130_fd_sc_hd__a21o_4
  _1643_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_31__.dout ),
    .B1(_0513_),
    .X(_0154_)
  );


  sky130_fd_sc_hd__and2_4
  _1644_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_32__.sout ),
    .X(_0514_)
  );


  sky130_fd_sc_hd__a21o_4
  _1645_
  (
    .A1(_0463_),
    .A2(mp[0]),
    .B1(_0514_),
    .X(\__BoundaryScanRegister_input_32__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1646_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_31__.sout ),
    .X(_0515_)
  );


  sky130_fd_sc_hd__a21o_4
  _1647_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_32__.dout ),
    .B1(_0515_),
    .X(_0155_)
  );


  sky130_fd_sc_hd__and2_4
  _1648_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_33__.sout ),
    .X(_0516_)
  );


  sky130_fd_sc_hd__a21o_4
  _1649_
  (
    .A1(_0463_),
    .A2(mp[1]),
    .B1(_0516_),
    .X(\__BoundaryScanRegister_input_33__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1650_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_32__.sout ),
    .X(_0517_)
  );


  sky130_fd_sc_hd__a21o_4
  _1651_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_33__.dout ),
    .B1(_0517_),
    .X(_0156_)
  );


  sky130_fd_sc_hd__and2_4
  _1652_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_34__.sout ),
    .X(_0518_)
  );


  sky130_fd_sc_hd__a21o_4
  _1653_
  (
    .A1(_0463_),
    .A2(mp[2]),
    .B1(_0518_),
    .X(\__BoundaryScanRegister_input_34__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1654_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_33__.sout ),
    .X(_0519_)
  );


  sky130_fd_sc_hd__a21o_4
  _1655_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_34__.dout ),
    .B1(_0519_),
    .X(_0157_)
  );


  sky130_fd_sc_hd__and2_4
  _1656_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_35__.sout ),
    .X(_0520_)
  );


  sky130_fd_sc_hd__a21o_4
  _1657_
  (
    .A1(_0463_),
    .A2(mp[3]),
    .B1(_0520_),
    .X(\__BoundaryScanRegister_input_35__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1658_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_34__.sout ),
    .X(_0521_)
  );


  sky130_fd_sc_hd__a21o_4
  _1659_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_35__.dout ),
    .B1(_0521_),
    .X(_0158_)
  );


  sky130_fd_sc_hd__and2_4
  _1660_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_36__.sout ),
    .X(_0522_)
  );


  sky130_fd_sc_hd__a21o_4
  _1661_
  (
    .A1(_0463_),
    .A2(mp[4]),
    .B1(_0522_),
    .X(\__BoundaryScanRegister_input_36__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1662_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_35__.sout ),
    .X(_0523_)
  );


  sky130_fd_sc_hd__a21o_4
  _1663_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_36__.dout ),
    .B1(_0523_),
    .X(_0159_)
  );


  sky130_fd_sc_hd__and2_4
  _1664_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_37__.sout ),
    .X(_0524_)
  );


  sky130_fd_sc_hd__a21o_4
  _1665_
  (
    .A1(_0463_),
    .A2(mp[5]),
    .B1(_0524_),
    .X(\__BoundaryScanRegister_input_37__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1666_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_36__.sout ),
    .X(_0525_)
  );


  sky130_fd_sc_hd__a21o_4
  _1667_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_37__.dout ),
    .B1(_0525_),
    .X(_0160_)
  );


  sky130_fd_sc_hd__and2_4
  _1668_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_38__.sout ),
    .X(_0526_)
  );


  sky130_fd_sc_hd__a21o_4
  _1669_
  (
    .A1(_0463_),
    .A2(mp[6]),
    .B1(_0526_),
    .X(\__BoundaryScanRegister_input_38__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1670_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_37__.sout ),
    .X(_0527_)
  );


  sky130_fd_sc_hd__a21o_4
  _1671_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_38__.dout ),
    .B1(_0527_),
    .X(_0161_)
  );


  sky130_fd_sc_hd__and2_4
  _1672_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_39__.sout ),
    .X(_0528_)
  );


  sky130_fd_sc_hd__a21o_4
  _1673_
  (
    .A1(_0463_),
    .A2(mp[7]),
    .B1(_0528_),
    .X(\__BoundaryScanRegister_input_39__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1674_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_38__.sout ),
    .X(_0529_)
  );


  sky130_fd_sc_hd__a21o_4
  _1675_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_39__.dout ),
    .B1(_0529_),
    .X(_0162_)
  );


  sky130_fd_sc_hd__and2_4
  _1676_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_3__.sout ),
    .X(_0530_)
  );


  sky130_fd_sc_hd__a21o_4
  _1677_
  (
    .A1(_0463_),
    .A2(mc[3]),
    .B1(_0530_),
    .X(\__BoundaryScanRegister_input_3__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1678_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_2__.sout ),
    .X(_0531_)
  );


  sky130_fd_sc_hd__a21o_4
  _1679_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_3__.dout ),
    .B1(_0531_),
    .X(_0163_)
  );


  sky130_fd_sc_hd__and2_4
  _1680_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_40__.sout ),
    .X(_0532_)
  );


  sky130_fd_sc_hd__a21o_4
  _1681_
  (
    .A1(_0463_),
    .A2(mp[8]),
    .B1(_0532_),
    .X(\__BoundaryScanRegister_input_40__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1682_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_39__.sout ),
    .X(_0533_)
  );


  sky130_fd_sc_hd__a21o_4
  _1683_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_40__.dout ),
    .B1(_0533_),
    .X(_0164_)
  );


  sky130_fd_sc_hd__and2_4
  _1684_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_41__.sout ),
    .X(_0534_)
  );


  sky130_fd_sc_hd__a21o_4
  _1685_
  (
    .A1(_0463_),
    .A2(mp[9]),
    .B1(_0534_),
    .X(\__BoundaryScanRegister_input_41__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1686_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_40__.sout ),
    .X(_0535_)
  );


  sky130_fd_sc_hd__a21o_4
  _1687_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_41__.dout ),
    .B1(_0535_),
    .X(_0165_)
  );


  sky130_fd_sc_hd__and2_4
  _1688_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_42__.sout ),
    .X(_0536_)
  );


  sky130_fd_sc_hd__a21o_4
  _1689_
  (
    .A1(_0463_),
    .A2(mp[10]),
    .B1(_0536_),
    .X(\__BoundaryScanRegister_input_42__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1690_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_41__.sout ),
    .X(_0537_)
  );


  sky130_fd_sc_hd__a21o_4
  _1691_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_42__.dout ),
    .B1(_0537_),
    .X(_0166_)
  );


  sky130_fd_sc_hd__and2_4
  _1692_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_43__.sout ),
    .X(_0538_)
  );


  sky130_fd_sc_hd__a21o_4
  _1693_
  (
    .A1(_0463_),
    .A2(mp[11]),
    .B1(_0538_),
    .X(\__BoundaryScanRegister_input_43__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1694_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_42__.sout ),
    .X(_0539_)
  );


  sky130_fd_sc_hd__a21o_4
  _1695_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_43__.dout ),
    .B1(_0539_),
    .X(_0167_)
  );


  sky130_fd_sc_hd__and2_4
  _1696_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_44__.sout ),
    .X(_0540_)
  );


  sky130_fd_sc_hd__a21o_4
  _1697_
  (
    .A1(_0463_),
    .A2(mp[12]),
    .B1(_0540_),
    .X(\__BoundaryScanRegister_input_44__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1698_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_43__.sout ),
    .X(_0541_)
  );


  sky130_fd_sc_hd__a21o_4
  _1699_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_44__.dout ),
    .B1(_0541_),
    .X(_0168_)
  );


  sky130_fd_sc_hd__and2_4
  _1700_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_45__.sout ),
    .X(_0542_)
  );


  sky130_fd_sc_hd__a21o_4
  _1701_
  (
    .A1(_0463_),
    .A2(mp[13]),
    .B1(_0542_),
    .X(\__BoundaryScanRegister_input_45__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1702_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_44__.sout ),
    .X(_0543_)
  );


  sky130_fd_sc_hd__a21o_4
  _1703_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_45__.dout ),
    .B1(_0543_),
    .X(_0169_)
  );


  sky130_fd_sc_hd__and2_4
  _1704_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_46__.sout ),
    .X(_0544_)
  );


  sky130_fd_sc_hd__a21o_4
  _1705_
  (
    .A1(_0463_),
    .A2(mp[14]),
    .B1(_0544_),
    .X(\__BoundaryScanRegister_input_46__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1706_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_45__.sout ),
    .X(_0545_)
  );


  sky130_fd_sc_hd__a21o_4
  _1707_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_46__.dout ),
    .B1(_0545_),
    .X(_0170_)
  );


  sky130_fd_sc_hd__and2_4
  _1708_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_47__.sout ),
    .X(_0546_)
  );


  sky130_fd_sc_hd__a21o_4
  _1709_
  (
    .A1(_0463_),
    .A2(mp[15]),
    .B1(_0546_),
    .X(\__BoundaryScanRegister_input_47__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1710_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_46__.sout ),
    .X(_0547_)
  );


  sky130_fd_sc_hd__a21o_4
  _1711_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_47__.dout ),
    .B1(_0547_),
    .X(_0171_)
  );


  sky130_fd_sc_hd__and2_4
  _1712_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_48__.sout ),
    .X(_0548_)
  );


  sky130_fd_sc_hd__a21o_4
  _1713_
  (
    .A1(_0463_),
    .A2(mp[16]),
    .B1(_0548_),
    .X(\__BoundaryScanRegister_input_48__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1714_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_47__.sout ),
    .X(_0549_)
  );


  sky130_fd_sc_hd__a21o_4
  _1715_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_48__.dout ),
    .B1(_0549_),
    .X(_0172_)
  );


  sky130_fd_sc_hd__and2_4
  _1716_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_49__.sout ),
    .X(_0550_)
  );


  sky130_fd_sc_hd__a21o_4
  _1717_
  (
    .A1(_0463_),
    .A2(mp[17]),
    .B1(_0550_),
    .X(\__BoundaryScanRegister_input_49__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1718_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_48__.sout ),
    .X(_0551_)
  );


  sky130_fd_sc_hd__a21o_4
  _1719_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_49__.dout ),
    .B1(_0551_),
    .X(_0173_)
  );


  sky130_fd_sc_hd__and2_4
  _1720_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_4__.sout ),
    .X(_0552_)
  );


  sky130_fd_sc_hd__a21o_4
  _1721_
  (
    .A1(_0463_),
    .A2(mc[4]),
    .B1(_0552_),
    .X(\__BoundaryScanRegister_input_4__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1722_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_3__.sout ),
    .X(_0553_)
  );


  sky130_fd_sc_hd__a21o_4
  _1723_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_4__.dout ),
    .B1(_0553_),
    .X(_0174_)
  );


  sky130_fd_sc_hd__and2_4
  _1724_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_50__.sout ),
    .X(_0554_)
  );


  sky130_fd_sc_hd__a21o_4
  _1725_
  (
    .A1(_0463_),
    .A2(mp[18]),
    .B1(_0554_),
    .X(\__BoundaryScanRegister_input_50__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1726_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_49__.sout ),
    .X(_0555_)
  );


  sky130_fd_sc_hd__a21o_4
  _1727_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_50__.dout ),
    .B1(_0555_),
    .X(_0175_)
  );


  sky130_fd_sc_hd__and2_4
  _1728_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_51__.sout ),
    .X(_0556_)
  );


  sky130_fd_sc_hd__a21o_4
  _1729_
  (
    .A1(_0463_),
    .A2(mp[19]),
    .B1(_0556_),
    .X(\__BoundaryScanRegister_input_51__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1730_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_50__.sout ),
    .X(_0557_)
  );


  sky130_fd_sc_hd__a21o_4
  _1731_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_51__.dout ),
    .B1(_0557_),
    .X(_0176_)
  );


  sky130_fd_sc_hd__and2_4
  _1732_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_52__.sout ),
    .X(_0558_)
  );


  sky130_fd_sc_hd__a21o_4
  _1733_
  (
    .A1(_0463_),
    .A2(mp[20]),
    .B1(_0558_),
    .X(\__BoundaryScanRegister_input_52__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1734_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_51__.sout ),
    .X(_0559_)
  );


  sky130_fd_sc_hd__a21o_4
  _1735_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_52__.dout ),
    .B1(_0559_),
    .X(_0177_)
  );


  sky130_fd_sc_hd__and2_4
  _1736_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_53__.sout ),
    .X(_0560_)
  );


  sky130_fd_sc_hd__a21o_4
  _1737_
  (
    .A1(_0463_),
    .A2(mp[21]),
    .B1(_0560_),
    .X(\__BoundaryScanRegister_input_53__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1738_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_52__.sout ),
    .X(_0561_)
  );


  sky130_fd_sc_hd__a21o_4
  _1739_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_53__.dout ),
    .B1(_0561_),
    .X(_0178_)
  );


  sky130_fd_sc_hd__and2_4
  _1740_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_54__.sout ),
    .X(_0562_)
  );


  sky130_fd_sc_hd__a21o_4
  _1741_
  (
    .A1(_0463_),
    .A2(mp[22]),
    .B1(_0562_),
    .X(\__BoundaryScanRegister_input_54__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1742_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_53__.sout ),
    .X(_0563_)
  );


  sky130_fd_sc_hd__a21o_4
  _1743_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_54__.dout ),
    .B1(_0563_),
    .X(_0179_)
  );


  sky130_fd_sc_hd__and2_4
  _1744_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_55__.sout ),
    .X(_0564_)
  );


  sky130_fd_sc_hd__a21o_4
  _1745_
  (
    .A1(_0463_),
    .A2(mp[23]),
    .B1(_0564_),
    .X(\__BoundaryScanRegister_input_55__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1746_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_54__.sout ),
    .X(_0565_)
  );


  sky130_fd_sc_hd__a21o_4
  _1747_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_55__.dout ),
    .B1(_0565_),
    .X(_0180_)
  );


  sky130_fd_sc_hd__and2_4
  _1748_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_56__.sout ),
    .X(_0566_)
  );


  sky130_fd_sc_hd__a21o_4
  _1749_
  (
    .A1(_0463_),
    .A2(mp[24]),
    .B1(_0566_),
    .X(\__BoundaryScanRegister_input_56__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1750_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_55__.sout ),
    .X(_0567_)
  );


  sky130_fd_sc_hd__a21o_4
  _1751_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_56__.dout ),
    .B1(_0567_),
    .X(_0181_)
  );


  sky130_fd_sc_hd__and2_4
  _1752_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_57__.sout ),
    .X(_0568_)
  );


  sky130_fd_sc_hd__a21o_4
  _1753_
  (
    .A1(_0463_),
    .A2(mp[25]),
    .B1(_0568_),
    .X(\__BoundaryScanRegister_input_57__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1754_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_56__.sout ),
    .X(_0569_)
  );


  sky130_fd_sc_hd__a21o_4
  _1755_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_57__.dout ),
    .B1(_0569_),
    .X(_0182_)
  );


  sky130_fd_sc_hd__and2_4
  _1756_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_58__.sout ),
    .X(_0570_)
  );


  sky130_fd_sc_hd__a21o_4
  _1757_
  (
    .A1(_0463_),
    .A2(mp[26]),
    .B1(_0570_),
    .X(\__BoundaryScanRegister_input_58__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1758_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_57__.sout ),
    .X(_0571_)
  );


  sky130_fd_sc_hd__a21o_4
  _1759_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_58__.dout ),
    .B1(_0571_),
    .X(_0183_)
  );


  sky130_fd_sc_hd__and2_4
  _1760_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_59__.sout ),
    .X(_0572_)
  );


  sky130_fd_sc_hd__a21o_4
  _1761_
  (
    .A1(_0463_),
    .A2(mp[27]),
    .B1(_0572_),
    .X(\__BoundaryScanRegister_input_59__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1762_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_58__.sout ),
    .X(_0573_)
  );


  sky130_fd_sc_hd__a21o_4
  _1763_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_59__.dout ),
    .B1(_0573_),
    .X(_0184_)
  );


  sky130_fd_sc_hd__and2_4
  _1764_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_5__.sout ),
    .X(_0574_)
  );


  sky130_fd_sc_hd__a21o_4
  _1765_
  (
    .A1(_0463_),
    .A2(mc[5]),
    .B1(_0574_),
    .X(\__BoundaryScanRegister_input_5__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1766_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_4__.sout ),
    .X(_0575_)
  );


  sky130_fd_sc_hd__a21o_4
  _1767_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_5__.dout ),
    .B1(_0575_),
    .X(_0185_)
  );


  sky130_fd_sc_hd__and2_4
  _1768_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_60__.sout ),
    .X(_0576_)
  );


  sky130_fd_sc_hd__a21o_4
  _1769_
  (
    .A1(_0463_),
    .A2(mp[28]),
    .B1(_0576_),
    .X(\__BoundaryScanRegister_input_60__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1770_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_59__.sout ),
    .X(_0577_)
  );


  sky130_fd_sc_hd__a21o_4
  _1771_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_60__.dout ),
    .B1(_0577_),
    .X(_0186_)
  );


  sky130_fd_sc_hd__and2_4
  _1772_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_61__.sout ),
    .X(_0578_)
  );


  sky130_fd_sc_hd__a21o_4
  _1773_
  (
    .A1(_0463_),
    .A2(mp[29]),
    .B1(_0578_),
    .X(\__BoundaryScanRegister_input_61__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1774_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_60__.sout ),
    .X(_0579_)
  );


  sky130_fd_sc_hd__a21o_4
  _1775_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_61__.dout ),
    .B1(_0579_),
    .X(_0187_)
  );


  sky130_fd_sc_hd__and2_4
  _1776_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_62__.sout ),
    .X(_0580_)
  );


  sky130_fd_sc_hd__a21o_4
  _1777_
  (
    .A1(_0463_),
    .A2(mp[30]),
    .B1(_0580_),
    .X(\__BoundaryScanRegister_input_62__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1778_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_61__.sout ),
    .X(_0581_)
  );


  sky130_fd_sc_hd__a21o_4
  _1779_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_62__.dout ),
    .B1(_0581_),
    .X(_0188_)
  );


  sky130_fd_sc_hd__and2_4
  _1780_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_63__.sout ),
    .X(_0582_)
  );


  sky130_fd_sc_hd__a21o_4
  _1781_
  (
    .A1(_0463_),
    .A2(mp[31]),
    .B1(_0582_),
    .X(\__BoundaryScanRegister_input_63__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1782_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_62__.sout ),
    .X(_0583_)
  );


  sky130_fd_sc_hd__a21o_4
  _1783_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_63__.dout ),
    .B1(_0583_),
    .X(_0189_)
  );


  sky130_fd_sc_hd__and2_4
  _1784_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_64__.sout ),
    .X(_0584_)
  );


  sky130_fd_sc_hd__a21o_4
  _1785_
  (
    .A1(_0463_),
    .A2(start),
    .B1(_0584_),
    .X(\__BoundaryScanRegister_input_64__.dout )
  );


  sky130_fd_sc_hd__and2_4
  _1786_
  (
    .A(shift),
    .B(\__BoundaryScanRegister_input_63__.sout ),
    .X(_0585_)
  );


  sky130_fd_sc_hd__a21o_4
  _1787_
  (
    .A1(_0462_),
    .A2(\__BoundaryScanRegister_input_64__.dout ),
    .B1(_0585_),
    .X(_0190_)
  );


  sky130_fd_sc_hd__and2_4
  _1788_
  (
    .A(test),
    .B(\__BoundaryScanRegister_input_6__.sout ),
    .X(_0586_)
  );


  sky130_fd_sc_hd__a21o_4
  _1789_
  (
    .A1(_0463_),
    .A2(mc[6]),
    .B1(_0586_),
    .X(\__BoundaryScanRegister_input_6__.dout )
  );


  sky130_fd_sc_hd__dfrtp_4
  _1790_
  (
    .CLK(tck),
    .D(_0130_),
    .Q(\__BoundaryScanRegister_input_0__.sout ),
    .RESET_B(_0000_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1791_
  (
    .CLK(tck),
    .D(_0131_),
    .Q(\__BoundaryScanRegister_input_10__.sout ),
    .RESET_B(_0001_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1792_
  (
    .CLK(tck),
    .D(_0132_),
    .Q(\__BoundaryScanRegister_input_11__.sout ),
    .RESET_B(_0002_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1793_
  (
    .CLK(tck),
    .D(_0133_),
    .Q(\__BoundaryScanRegister_input_12__.sout ),
    .RESET_B(_0003_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1794_
  (
    .CLK(tck),
    .D(_0134_),
    .Q(\__BoundaryScanRegister_input_13__.sout ),
    .RESET_B(_0004_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1795_
  (
    .CLK(tck),
    .D(_0135_),
    .Q(\__BoundaryScanRegister_input_14__.sout ),
    .RESET_B(_0005_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1796_
  (
    .CLK(tck),
    .D(_0136_),
    .Q(\__BoundaryScanRegister_input_15__.sout ),
    .RESET_B(_0006_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1797_
  (
    .CLK(tck),
    .D(_0137_),
    .Q(\__BoundaryScanRegister_input_16__.sout ),
    .RESET_B(_0007_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1798_
  (
    .CLK(tck),
    .D(_0138_),
    .Q(\__BoundaryScanRegister_input_17__.sout ),
    .RESET_B(_0008_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1799_
  (
    .CLK(tck),
    .D(_0139_),
    .Q(\__BoundaryScanRegister_input_18__.sout ),
    .RESET_B(_0009_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1800_
  (
    .CLK(tck),
    .D(_0140_),
    .Q(\__BoundaryScanRegister_input_19__.sout ),
    .RESET_B(_0010_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1801_
  (
    .CLK(tck),
    .D(_0141_),
    .Q(\__BoundaryScanRegister_input_1__.sout ),
    .RESET_B(_0011_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1802_
  (
    .CLK(tck),
    .D(_0142_),
    .Q(\__BoundaryScanRegister_input_20__.sout ),
    .RESET_B(_0012_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1803_
  (
    .CLK(tck),
    .D(_0143_),
    .Q(\__BoundaryScanRegister_input_21__.sout ),
    .RESET_B(_0013_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1804_
  (
    .CLK(tck),
    .D(_0144_),
    .Q(\__BoundaryScanRegister_input_22__.sout ),
    .RESET_B(_0014_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1805_
  (
    .CLK(tck),
    .D(_0145_),
    .Q(\__BoundaryScanRegister_input_23__.sout ),
    .RESET_B(_0015_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1806_
  (
    .CLK(tck),
    .D(_0146_),
    .Q(\__BoundaryScanRegister_input_24__.sout ),
    .RESET_B(_0016_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1807_
  (
    .CLK(tck),
    .D(_0147_),
    .Q(\__BoundaryScanRegister_input_25__.sout ),
    .RESET_B(_0017_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1808_
  (
    .CLK(tck),
    .D(_0148_),
    .Q(\__BoundaryScanRegister_input_26__.sout ),
    .RESET_B(_0018_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1809_
  (
    .CLK(tck),
    .D(_0149_),
    .Q(\__BoundaryScanRegister_input_27__.sout ),
    .RESET_B(_0019_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1810_
  (
    .CLK(tck),
    .D(_0150_),
    .Q(\__BoundaryScanRegister_input_28__.sout ),
    .RESET_B(_0020_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1811_
  (
    .CLK(tck),
    .D(_0151_),
    .Q(\__BoundaryScanRegister_input_29__.sout ),
    .RESET_B(_0021_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1812_
  (
    .CLK(tck),
    .D(_0152_),
    .Q(\__BoundaryScanRegister_input_2__.sout ),
    .RESET_B(_0022_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1813_
  (
    .CLK(tck),
    .D(_0153_),
    .Q(\__BoundaryScanRegister_input_30__.sout ),
    .RESET_B(_0023_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1814_
  (
    .CLK(tck),
    .D(_0154_),
    .Q(\__BoundaryScanRegister_input_31__.sout ),
    .RESET_B(_0024_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1815_
  (
    .CLK(tck),
    .D(_0155_),
    .Q(\__BoundaryScanRegister_input_32__.sout ),
    .RESET_B(_0025_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1816_
  (
    .CLK(tck),
    .D(_0156_),
    .Q(\__BoundaryScanRegister_input_33__.sout ),
    .RESET_B(_0026_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1817_
  (
    .CLK(tck),
    .D(_0157_),
    .Q(\__BoundaryScanRegister_input_34__.sout ),
    .RESET_B(_0027_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1818_
  (
    .CLK(tck),
    .D(_0158_),
    .Q(\__BoundaryScanRegister_input_35__.sout ),
    .RESET_B(_0028_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1819_
  (
    .CLK(tck),
    .D(_0159_),
    .Q(\__BoundaryScanRegister_input_36__.sout ),
    .RESET_B(_0029_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1820_
  (
    .CLK(tck),
    .D(_0160_),
    .Q(\__BoundaryScanRegister_input_37__.sout ),
    .RESET_B(_0030_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1821_
  (
    .CLK(tck),
    .D(_0161_),
    .Q(\__BoundaryScanRegister_input_38__.sout ),
    .RESET_B(_0031_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1822_
  (
    .CLK(tck),
    .D(_0162_),
    .Q(\__BoundaryScanRegister_input_39__.sout ),
    .RESET_B(_0032_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1823_
  (
    .CLK(tck),
    .D(_0163_),
    .Q(\__BoundaryScanRegister_input_3__.sout ),
    .RESET_B(_0033_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1824_
  (
    .CLK(tck),
    .D(_0164_),
    .Q(\__BoundaryScanRegister_input_40__.sout ),
    .RESET_B(_0034_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1825_
  (
    .CLK(tck),
    .D(_0165_),
    .Q(\__BoundaryScanRegister_input_41__.sout ),
    .RESET_B(_0035_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1826_
  (
    .CLK(tck),
    .D(_0166_),
    .Q(\__BoundaryScanRegister_input_42__.sout ),
    .RESET_B(_0036_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1827_
  (
    .CLK(tck),
    .D(_0167_),
    .Q(\__BoundaryScanRegister_input_43__.sout ),
    .RESET_B(_0037_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1828_
  (
    .CLK(tck),
    .D(_0168_),
    .Q(\__BoundaryScanRegister_input_44__.sout ),
    .RESET_B(_0038_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1829_
  (
    .CLK(tck),
    .D(_0169_),
    .Q(\__BoundaryScanRegister_input_45__.sout ),
    .RESET_B(_0039_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1830_
  (
    .CLK(tck),
    .D(_0170_),
    .Q(\__BoundaryScanRegister_input_46__.sout ),
    .RESET_B(_0040_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1831_
  (
    .CLK(tck),
    .D(_0171_),
    .Q(\__BoundaryScanRegister_input_47__.sout ),
    .RESET_B(_0041_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1832_
  (
    .CLK(tck),
    .D(_0172_),
    .Q(\__BoundaryScanRegister_input_48__.sout ),
    .RESET_B(_0042_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1833_
  (
    .CLK(tck),
    .D(_0173_),
    .Q(\__BoundaryScanRegister_input_49__.sout ),
    .RESET_B(_0043_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1834_
  (
    .CLK(tck),
    .D(_0174_),
    .Q(\__BoundaryScanRegister_input_4__.sout ),
    .RESET_B(_0044_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1835_
  (
    .CLK(tck),
    .D(_0175_),
    .Q(\__BoundaryScanRegister_input_50__.sout ),
    .RESET_B(_0045_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1836_
  (
    .CLK(tck),
    .D(_0176_),
    .Q(\__BoundaryScanRegister_input_51__.sout ),
    .RESET_B(_0046_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1837_
  (
    .CLK(tck),
    .D(_0177_),
    .Q(\__BoundaryScanRegister_input_52__.sout ),
    .RESET_B(_0047_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1838_
  (
    .CLK(tck),
    .D(_0178_),
    .Q(\__BoundaryScanRegister_input_53__.sout ),
    .RESET_B(_0048_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1839_
  (
    .CLK(tck),
    .D(_0179_),
    .Q(\__BoundaryScanRegister_input_54__.sout ),
    .RESET_B(_0049_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1840_
  (
    .CLK(tck),
    .D(_0180_),
    .Q(\__BoundaryScanRegister_input_55__.sout ),
    .RESET_B(_0050_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1841_
  (
    .CLK(tck),
    .D(_0181_),
    .Q(\__BoundaryScanRegister_input_56__.sout ),
    .RESET_B(_0051_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1842_
  (
    .CLK(tck),
    .D(_0182_),
    .Q(\__BoundaryScanRegister_input_57__.sout ),
    .RESET_B(_0052_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1843_
  (
    .CLK(tck),
    .D(_0183_),
    .Q(\__BoundaryScanRegister_input_58__.sout ),
    .RESET_B(_0053_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1844_
  (
    .CLK(tck),
    .D(_0184_),
    .Q(\__BoundaryScanRegister_input_59__.sout ),
    .RESET_B(_0054_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1845_
  (
    .CLK(tck),
    .D(_0185_),
    .Q(\__BoundaryScanRegister_input_5__.sout ),
    .RESET_B(_0055_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1846_
  (
    .CLK(tck),
    .D(_0186_),
    .Q(\__BoundaryScanRegister_input_60__.sout ),
    .RESET_B(_0056_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1847_
  (
    .CLK(tck),
    .D(_0187_),
    .Q(\__BoundaryScanRegister_input_61__.sout ),
    .RESET_B(_0057_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1848_
  (
    .CLK(tck),
    .D(_0188_),
    .Q(\__BoundaryScanRegister_input_62__.sout ),
    .RESET_B(_0058_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1849_
  (
    .CLK(tck),
    .D(_0189_),
    .Q(\__BoundaryScanRegister_input_63__.sout ),
    .RESET_B(_0059_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1850_
  (
    .CLK(tck),
    .D(_0190_),
    .Q(\__BoundaryScanRegister_input_64__.sout ),
    .RESET_B(_0060_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1851_
  (
    .CLK(tck),
    .D(_0191_),
    .Q(\__BoundaryScanRegister_input_6__.sout ),
    .RESET_B(_0061_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1852_
  (
    .CLK(tck),
    .D(_0192_),
    .Q(\__BoundaryScanRegister_input_7__.sout ),
    .RESET_B(_0062_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1853_
  (
    .CLK(tck),
    .D(_0193_),
    .Q(\__BoundaryScanRegister_input_8__.sout ),
    .RESET_B(_0063_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1854_
  (
    .CLK(tck),
    .D(_0194_),
    .Q(\__BoundaryScanRegister_input_10__.sin ),
    .RESET_B(_0064_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1855_
  (
    .CLK(tck),
    .D(_0195_),
    .Q(\__BoundaryScanRegister_output_100__.sout ),
    .RESET_B(_0065_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1856_
  (
    .CLK(tck),
    .D(_0196_),
    .Q(\__BoundaryScanRegister_output_101__.sout ),
    .RESET_B(_0066_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1857_
  (
    .CLK(tck),
    .D(_0197_),
    .Q(\__BoundaryScanRegister_output_102__.sout ),
    .RESET_B(_0067_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1858_
  (
    .CLK(tck),
    .D(_0198_),
    .Q(\__BoundaryScanRegister_output_103__.sout ),
    .RESET_B(_0068_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1859_
  (
    .CLK(tck),
    .D(_0199_),
    .Q(\__BoundaryScanRegister_output_104__.sout ),
    .RESET_B(_0069_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1860_
  (
    .CLK(tck),
    .D(_0200_),
    .Q(\__BoundaryScanRegister_output_105__.sout ),
    .RESET_B(_0070_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1861_
  (
    .CLK(tck),
    .D(_0201_),
    .Q(\__BoundaryScanRegister_output_106__.sout ),
    .RESET_B(_0071_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1862_
  (
    .CLK(tck),
    .D(_0202_),
    .Q(\__BoundaryScanRegister_output_107__.sout ),
    .RESET_B(_0072_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1863_
  (
    .CLK(tck),
    .D(_0203_),
    .Q(\__BoundaryScanRegister_output_108__.sout ),
    .RESET_B(_0073_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1864_
  (
    .CLK(tck),
    .D(_0204_),
    .Q(\__BoundaryScanRegister_output_109__.sout ),
    .RESET_B(_0074_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1865_
  (
    .CLK(tck),
    .D(_0205_),
    .Q(\__BoundaryScanRegister_output_110__.sout ),
    .RESET_B(_0075_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1866_
  (
    .CLK(tck),
    .D(_0206_),
    .Q(\__BoundaryScanRegister_output_111__.sout ),
    .RESET_B(_0076_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1867_
  (
    .CLK(tck),
    .D(_0207_),
    .Q(\__BoundaryScanRegister_output_112__.sout ),
    .RESET_B(_0077_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1868_
  (
    .CLK(tck),
    .D(_0208_),
    .Q(\__BoundaryScanRegister_output_113__.sout ),
    .RESET_B(_0078_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1869_
  (
    .CLK(tck),
    .D(_0209_),
    .Q(\__BoundaryScanRegister_output_114__.sout ),
    .RESET_B(_0079_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1870_
  (
    .CLK(tck),
    .D(_0210_),
    .Q(\__BoundaryScanRegister_output_115__.sout ),
    .RESET_B(_0080_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1871_
  (
    .CLK(tck),
    .D(_0211_),
    .Q(\__BoundaryScanRegister_output_116__.sout ),
    .RESET_B(_0081_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1872_
  (
    .CLK(tck),
    .D(_0212_),
    .Q(\__BoundaryScanRegister_output_117__.sout ),
    .RESET_B(_0082_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1873_
  (
    .CLK(tck),
    .D(_0213_),
    .Q(\__BoundaryScanRegister_output_118__.sout ),
    .RESET_B(_0083_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1874_
  (
    .CLK(tck),
    .D(_0214_),
    .Q(\__BoundaryScanRegister_output_119__.sout ),
    .RESET_B(_0084_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1875_
  (
    .CLK(tck),
    .D(_0215_),
    .Q(\__BoundaryScanRegister_output_120__.sout ),
    .RESET_B(_0085_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1876_
  (
    .CLK(tck),
    .D(_0216_),
    .Q(\__BoundaryScanRegister_output_121__.sout ),
    .RESET_B(_0086_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1877_
  (
    .CLK(tck),
    .D(_0217_),
    .Q(\__BoundaryScanRegister_output_122__.sout ),
    .RESET_B(_0087_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1878_
  (
    .CLK(tck),
    .D(_0218_),
    .Q(\__BoundaryScanRegister_output_123__.sout ),
    .RESET_B(_0088_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1879_
  (
    .CLK(tck),
    .D(_0219_),
    .Q(\__BoundaryScanRegister_output_124__.sout ),
    .RESET_B(_0089_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1880_
  (
    .CLK(tck),
    .D(_0220_),
    .Q(\__BoundaryScanRegister_output_125__.sout ),
    .RESET_B(_0090_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1881_
  (
    .CLK(tck),
    .D(_0221_),
    .Q(\__BoundaryScanRegister_output_126__.sout ),
    .RESET_B(_0091_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1882_
  (
    .CLK(tck),
    .D(_0222_),
    .Q(\__BoundaryScanRegister_output_127__.sout ),
    .RESET_B(_0092_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1883_
  (
    .CLK(tck),
    .D(_0223_),
    .Q(\__BoundaryScanRegister_output_128__.sout ),
    .RESET_B(_0093_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1884_
  (
    .CLK(tck),
    .D(_0224_),
    .Q(sout),
    .RESET_B(_0094_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1885_
  (
    .CLK(tck),
    .D(_0225_),
    .Q(\__BoundaryScanRegister_output_65__.sout ),
    .RESET_B(_0095_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1886_
  (
    .CLK(tck),
    .D(_0226_),
    .Q(\__BoundaryScanRegister_output_66__.sout ),
    .RESET_B(_0096_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1887_
  (
    .CLK(tck),
    .D(_0227_),
    .Q(\__BoundaryScanRegister_output_67__.sout ),
    .RESET_B(_0097_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1888_
  (
    .CLK(tck),
    .D(_0228_),
    .Q(\__BoundaryScanRegister_output_68__.sout ),
    .RESET_B(_0098_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1889_
  (
    .CLK(tck),
    .D(_0229_),
    .Q(\__BoundaryScanRegister_output_69__.sout ),
    .RESET_B(_0099_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1890_
  (
    .CLK(tck),
    .D(_0230_),
    .Q(\__BoundaryScanRegister_output_70__.sout ),
    .RESET_B(_0100_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1891_
  (
    .CLK(tck),
    .D(_0231_),
    .Q(\__BoundaryScanRegister_output_71__.sout ),
    .RESET_B(_0101_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1892_
  (
    .CLK(tck),
    .D(_0232_),
    .Q(\__BoundaryScanRegister_output_72__.sout ),
    .RESET_B(_0102_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1893_
  (
    .CLK(tck),
    .D(_0233_),
    .Q(\__BoundaryScanRegister_output_73__.sout ),
    .RESET_B(_0103_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1894_
  (
    .CLK(tck),
    .D(_0234_),
    .Q(\__BoundaryScanRegister_output_74__.sout ),
    .RESET_B(_0104_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1895_
  (
    .CLK(tck),
    .D(_0235_),
    .Q(\__BoundaryScanRegister_output_75__.sout ),
    .RESET_B(_0105_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1896_
  (
    .CLK(tck),
    .D(_0236_),
    .Q(\__BoundaryScanRegister_output_76__.sout ),
    .RESET_B(_0106_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1897_
  (
    .CLK(tck),
    .D(_0237_),
    .Q(\__BoundaryScanRegister_output_77__.sout ),
    .RESET_B(_0107_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1898_
  (
    .CLK(tck),
    .D(_0238_),
    .Q(\__BoundaryScanRegister_output_78__.sout ),
    .RESET_B(_0108_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1899_
  (
    .CLK(tck),
    .D(_0239_),
    .Q(\__BoundaryScanRegister_output_79__.sout ),
    .RESET_B(_0109_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1900_
  (
    .CLK(tck),
    .D(_0240_),
    .Q(\__BoundaryScanRegister_output_80__.sout ),
    .RESET_B(_0110_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1901_
  (
    .CLK(tck),
    .D(_0241_),
    .Q(\__BoundaryScanRegister_output_81__.sout ),
    .RESET_B(_0111_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1902_
  (
    .CLK(tck),
    .D(_0242_),
    .Q(\__BoundaryScanRegister_output_82__.sout ),
    .RESET_B(_0112_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1903_
  (
    .CLK(tck),
    .D(_0243_),
    .Q(\__BoundaryScanRegister_output_83__.sout ),
    .RESET_B(_0113_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1904_
  (
    .CLK(tck),
    .D(_0244_),
    .Q(\__BoundaryScanRegister_output_84__.sout ),
    .RESET_B(_0114_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1905_
  (
    .CLK(tck),
    .D(_0245_),
    .Q(\__BoundaryScanRegister_output_85__.sout ),
    .RESET_B(_0115_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1906_
  (
    .CLK(tck),
    .D(_0246_),
    .Q(\__BoundaryScanRegister_output_86__.sout ),
    .RESET_B(_0116_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1907_
  (
    .CLK(tck),
    .D(_0247_),
    .Q(\__BoundaryScanRegister_output_87__.sout ),
    .RESET_B(_0117_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1908_
  (
    .CLK(tck),
    .D(_0248_),
    .Q(\__BoundaryScanRegister_output_88__.sout ),
    .RESET_B(_0118_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1909_
  (
    .CLK(tck),
    .D(_0249_),
    .Q(\__BoundaryScanRegister_output_89__.sout ),
    .RESET_B(_0119_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1910_
  (
    .CLK(tck),
    .D(_0250_),
    .Q(\__BoundaryScanRegister_output_90__.sout ),
    .RESET_B(_0120_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1911_
  (
    .CLK(tck),
    .D(_0251_),
    .Q(\__BoundaryScanRegister_output_91__.sout ),
    .RESET_B(_0121_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1912_
  (
    .CLK(tck),
    .D(_0252_),
    .Q(\__BoundaryScanRegister_output_92__.sout ),
    .RESET_B(_0122_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1913_
  (
    .CLK(tck),
    .D(_0253_),
    .Q(\__BoundaryScanRegister_output_93__.sout ),
    .RESET_B(_0123_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1914_
  (
    .CLK(tck),
    .D(_0254_),
    .Q(\__BoundaryScanRegister_output_94__.sout ),
    .RESET_B(_0124_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1915_
  (
    .CLK(tck),
    .D(_0255_),
    .Q(\__BoundaryScanRegister_output_95__.sout ),
    .RESET_B(_0125_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1916_
  (
    .CLK(tck),
    .D(_0256_),
    .Q(\__BoundaryScanRegister_output_96__.sout ),
    .RESET_B(_0126_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1917_
  (
    .CLK(tck),
    .D(_0257_),
    .Q(\__BoundaryScanRegister_output_97__.sout ),
    .RESET_B(_0127_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1918_
  (
    .CLK(tck),
    .D(_0258_),
    .Q(\__BoundaryScanRegister_output_98__.sout ),
    .RESET_B(_0128_)
  );


  sky130_fd_sc_hd__dfrtp_4
  _1919_
  (
    .CLK(tck),
    .D(_0259_),
    .Q(\__BoundaryScanRegister_output_100__.sin ),
    .RESET_B(_0129_)
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0882_ 
  (
    .A(\__uuf__.fsm.state[0] ),
    .Y(\__uuf__._0766_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0883_ 
  (
    .A(\__uuf__.count[1] ),
    .Y(\__uuf__._0767_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0884_ 
  (
    .A(\__BoundaryScanRegister_output_65__.sin ),
    .Y(\__uuf__._0768_ )
  );


  sky130_fd_sc_hd__or4_4
  \__uuf__._0885_ 
  (
    .A(\__uuf__._0768_ ),
    .B(\__uuf__.count[5] ),
    .C(\__uuf__.count[4] ),
    .D(\__uuf__.count[3] ),
    .X(\__uuf__._0769_ )
  );


  sky130_fd_sc_hd__or4_4
  \__uuf__._0886_ 
  (
    .A(\__uuf__.count[2] ),
    .B(\__uuf__._0767_ ),
    .C(\__uuf__.count[0] ),
    .D(\__uuf__._0769_ ),
    .X(\__uuf__._0770_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0887_ 
  (
    .A(\__uuf__._0770_ ),
    .Y(\__uuf__._0771_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._0888_ 
  (
    .A(\__uuf__._0766_ ),
    .B(\__uuf__.fsm.state[1] ),
    .C(\__uuf__._0771_ ),
    .X(\__uuf__._0772_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0889_ 
  (
    .A(\__uuf__._0772_ ),
    .Y(\__uuf__._0773_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0890_ 
  (
    .A(\__uuf__._0773_ ),
    .X(\__uuf__._0774_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0891_ 
  (
    .A(\__uuf__._0774_ ),
    .X(\__uuf__._0775_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0892_ 
  (
    .A(\__uuf__.count[2] ),
    .Y(\__uuf__._0776_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0893_ 
  (
    .A(\__uuf__.count[0] ),
    .Y(\__uuf__._0777_ )
  );


  sky130_fd_sc_hd__or2_4
  \__uuf__._0894_ 
  (
    .A(\__uuf__._0767_ ),
    .B(\__uuf__._0777_ ),
    .X(\__uuf__._0778_ )
  );


  sky130_fd_sc_hd__or2_4
  \__uuf__._0895_ 
  (
    .A(\__uuf__._0776_ ),
    .B(\__uuf__._0778_ ),
    .X(\__uuf__._0779_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0896_ 
  (
    .A(\__uuf__._0779_ ),
    .Y(\__uuf__._0780_ )
  );


  sky130_fd_sc_hd__and2_4
  \__uuf__._0897_ 
  (
    .A(\__uuf__.count[3] ),
    .B(\__uuf__._0780_ ),
    .X(\__uuf__._0781_ )
  );


  sky130_fd_sc_hd__and2_4
  \__uuf__._0898_ 
  (
    .A(\__uuf__.count[4] ),
    .B(\__uuf__._0781_ ),
    .X(\__uuf__._0782_ )
  );


  sky130_fd_sc_hd__and2_4
  \__uuf__._0899_ 
  (
    .A(\__uuf__.count[5] ),
    .B(\__uuf__._0782_ ),
    .X(\__uuf__._0783_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0900_ 
  (
    .A(\__uuf__._0783_ ),
    .Y(\__uuf__._0784_ )
  );


  sky130_fd_sc_hd__or2_4
  \__uuf__._0901_ 
  (
    .A(\__uuf__._0768_ ),
    .B(\__uuf__._0784_ ),
    .X(\__uuf__._0785_ )
  );


  sky130_fd_sc_hd__or2_4
  \__uuf__._0902_ 
  (
    .A(\__BoundaryScanRegister_output_65__.sin ),
    .B(\__uuf__._0783_ ),
    .X(\__uuf__._0786_ )
  );


  sky130_fd_sc_hd__or2_4
  \__uuf__._0903_ 
  (
    .A(\__uuf__.fsm.state[0] ),
    .B(\__uuf__.fsm.state[1] ),
    .X(\__uuf__._0787_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0904_ 
  (
    .A(\__uuf__._0787_ ),
    .Y(\__uuf__._0788_ )
  );


  sky130_fd_sc_hd__or2_4
  \__uuf__._0905_ 
  (
    .A(\__uuf__._0773_ ),
    .B(\__uuf__._0788_ ),
    .X(\__uuf__._0789_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0906_ 
  (
    .A(\__uuf__._0789_ ),
    .Y(\__uuf__._0790_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0907_ 
  (
    .A(\__uuf__._0790_ ),
    .X(\__uuf__._0791_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0908_ 
  (
    .A1(\__uuf__._0775_ ),
    .A2(\__uuf__._0785_ ),
    .A3(\__uuf__._0786_ ),
    .B1(\__BoundaryScanRegister_output_65__.sin ),
    .B2(\__uuf__._0791_ ),
    .X(\__uuf__._0431_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0909_ 
  (
    .A(rst),
    .Y(\__uuf__._0792_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0910_ 
  (
    .A(\__uuf__._0792_ ),
    .X(\__uuf__._0793_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0911_ 
  (
    .A(\__uuf__._0793_ ),
    .X(\__uuf__._0794_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0912_ 
  (
    .A(\__uuf__._0794_ ),
    .X(\__uuf__._0359_ )
  );


  sky130_fd_sc_hd__or2_4
  \__uuf__._0913_ 
  (
    .A(\__uuf__.count[5] ),
    .B(\__uuf__._0782_ ),
    .X(\__uuf__._0795_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0914_ 
  (
    .A1(\__uuf__._0774_ ),
    .A2(\__uuf__._0795_ ),
    .A3(\__uuf__._0784_ ),
    .B1(\__uuf__.count[5] ),
    .B2(\__uuf__._0791_ ),
    .X(\__uuf__._0430_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0915_ 
  (
    .A(\__uuf__._0359_ ),
    .X(\__uuf__._0358_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0916_ 
  (
    .A(\__uuf__._0782_ ),
    .Y(\__uuf__._0796_ )
  );


  sky130_fd_sc_hd__or2_4
  \__uuf__._0917_ 
  (
    .A(\__uuf__.count[4] ),
    .B(\__uuf__._0781_ ),
    .X(\__uuf__._0797_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0918_ 
  (
    .A1(\__uuf__._0796_ ),
    .A2(\__uuf__._0797_ ),
    .A3(\__uuf__._0775_ ),
    .B1(\__uuf__.count[4] ),
    .B2(\__uuf__._0791_ ),
    .X(\__uuf__._0429_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0919_ 
  (
    .A(\__uuf__._0359_ ),
    .X(\__uuf__._0357_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._0920_ 
  (
    .A(\__uuf__._0781_ ),
    .Y(\__uuf__._0798_ )
  );


  sky130_fd_sc_hd__or2_4
  \__uuf__._0921_ 
  (
    .A(\__uuf__.count[3] ),
    .B(\__uuf__._0780_ ),
    .X(\__uuf__._0799_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0922_ 
  (
    .A1(\__uuf__._0798_ ),
    .A2(\__uuf__._0799_ ),
    .A3(\__uuf__._0775_ ),
    .B1(\__uuf__.count[3] ),
    .B2(\__uuf__._0791_ ),
    .X(\__uuf__._0428_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0923_ 
  (
    .A(\__uuf__._0359_ ),
    .X(\__uuf__._0356_ )
  );


  sky130_fd_sc_hd__nand2_4
  \__uuf__._0924_ 
  (
    .A(\__uuf__._0776_ ),
    .B(\__uuf__._0778_ ),
    .Y(\__uuf__._0800_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0925_ 
  (
    .A1(\__uuf__._0779_ ),
    .A2(\__uuf__._0800_ ),
    .A3(\__uuf__._0775_ ),
    .B1(\__uuf__.count[2] ),
    .B2(\__uuf__._0790_ ),
    .X(\__uuf__._0427_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0926_ 
  (
    .A(\__uuf__._0359_ ),
    .X(\__uuf__._0355_ )
  );


  sky130_fd_sc_hd__or2_4
  \__uuf__._0927_ 
  (
    .A(\__uuf__.count[1] ),
    .B(\__uuf__.count[0] ),
    .X(\__uuf__._0801_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0928_ 
  (
    .A1(\__uuf__._0778_ ),
    .A2(\__uuf__._0801_ ),
    .A3(\__uuf__._0775_ ),
    .B1(\__uuf__.count[1] ),
    .B2(\__uuf__._0790_ ),
    .X(\__uuf__._0426_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0929_ 
  (
    .A(\__uuf__._0794_ ),
    .X(\__uuf__._0802_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0930_ 
  (
    .A(\__uuf__._0802_ ),
    .X(\__uuf__._0354_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0931_ 
  (
    .A(\__uuf__._0773_ ),
    .X(\__uuf__._0803_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0932_ 
  (
    .A(\__uuf__._0803_ ),
    .X(\__uuf__._0804_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._0933_ 
  (
    .A1(\__uuf__.count[0] ),
    .A2(\__uuf__._0804_ ),
    .B1(\__uuf__._0777_ ),
    .B2(\__uuf__._0791_ ),
    .X(\__uuf__._0425_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0934_ 
  (
    .A(\__uuf__._0802_ ),
    .X(\__uuf__._0353_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0935_ 
  (
    .A(\__uuf__._0772_ ),
    .X(\__uuf__._0805_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0936_ 
  (
    .A(\__uuf__._0805_ ),
    .X(\__uuf__._0806_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0937_ 
  (
    .A(\__uuf__._0787_ ),
    .X(\__uuf__._0807_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0938_ 
  (
    .A(\__uuf__._0807_ ),
    .X(\__uuf__._0808_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0939_ 
  (
    .A1(\__uuf__._0806_ ),
    .A2(\__uuf__._0808_ ),
    .A3(prod[63]),
    .B1(\__uuf__.multiplier.csa0.sum ),
    .B2(\__uuf__._0804_ ),
    .X(\__uuf__._0424_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0940_ 
  (
    .A(\__uuf__._0802_ ),
    .X(\__uuf__._0352_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0941_ 
  (
    .A1(\__uuf__._0806_ ),
    .A2(\__uuf__._0808_ ),
    .A3(prod[62]),
    .B1(prod[63]),
    .B2(\__uuf__._0804_ ),
    .X(\__uuf__._0423_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0942_ 
  (
    .A(\__uuf__._0802_ ),
    .X(\__uuf__._0351_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0943_ 
  (
    .A1(\__uuf__._0806_ ),
    .A2(\__uuf__._0808_ ),
    .A3(prod[61]),
    .B1(prod[62]),
    .B2(\__uuf__._0804_ ),
    .X(\__uuf__._0422_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0944_ 
  (
    .A(\__uuf__._0802_ ),
    .X(\__uuf__._0350_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0945_ 
  (
    .A1(\__uuf__._0806_ ),
    .A2(\__uuf__._0808_ ),
    .A3(prod[60]),
    .B1(prod[61]),
    .B2(\__uuf__._0804_ ),
    .X(\__uuf__._0421_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0946_ 
  (
    .A(\__uuf__._0794_ ),
    .X(\__uuf__._0809_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0947_ 
  (
    .A(\__uuf__._0809_ ),
    .X(\__uuf__._0349_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0948_ 
  (
    .A(\__uuf__._0774_ ),
    .X(\__uuf__._0810_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0949_ 
  (
    .A1(\__uuf__._0806_ ),
    .A2(\__uuf__._0808_ ),
    .A3(prod[59]),
    .B1(prod[60]),
    .B2(\__uuf__._0810_ ),
    .X(\__uuf__._0420_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0950_ 
  (
    .A(\__uuf__._0809_ ),
    .X(\__uuf__._0348_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0951_ 
  (
    .A(\__uuf__._0772_ ),
    .X(\__uuf__._0811_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0952_ 
  (
    .A(\__uuf__._0811_ ),
    .X(\__uuf__._0812_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0953_ 
  (
    .A(\__uuf__._0787_ ),
    .X(\__uuf__._0813_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0954_ 
  (
    .A(\__uuf__._0813_ ),
    .X(\__uuf__._0814_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0955_ 
  (
    .A1(\__uuf__._0812_ ),
    .A2(\__uuf__._0814_ ),
    .A3(prod[58]),
    .B1(prod[59]),
    .B2(\__uuf__._0810_ ),
    .X(\__uuf__._0419_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0956_ 
  (
    .A(\__uuf__._0809_ ),
    .X(\__uuf__._0347_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0957_ 
  (
    .A1(\__uuf__._0812_ ),
    .A2(\__uuf__._0814_ ),
    .A3(prod[57]),
    .B1(prod[58]),
    .B2(\__uuf__._0810_ ),
    .X(\__uuf__._0418_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0958_ 
  (
    .A(\__uuf__._0809_ ),
    .X(\__uuf__._0346_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0959_ 
  (
    .A1(\__uuf__._0812_ ),
    .A2(\__uuf__._0814_ ),
    .A3(prod[56]),
    .B1(prod[57]),
    .B2(\__uuf__._0810_ ),
    .X(\__uuf__._0417_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0960_ 
  (
    .A(\__uuf__._0809_ ),
    .X(\__uuf__._0345_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0961_ 
  (
    .A1(\__uuf__._0812_ ),
    .A2(\__uuf__._0814_ ),
    .A3(prod[55]),
    .B1(prod[56]),
    .B2(\__uuf__._0810_ ),
    .X(\__uuf__._0416_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0962_ 
  (
    .A(\__uuf__._0792_ ),
    .X(\__uuf__._0815_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0963_ 
  (
    .A(\__uuf__._0815_ ),
    .X(\__uuf__._0816_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0964_ 
  (
    .A(\__uuf__._0816_ ),
    .X(\__uuf__._0817_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0965_ 
  (
    .A(\__uuf__._0817_ ),
    .X(\__uuf__._0344_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0966_ 
  (
    .A(\__uuf__._0774_ ),
    .X(\__uuf__._0818_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0967_ 
  (
    .A1(\__uuf__._0812_ ),
    .A2(\__uuf__._0814_ ),
    .A3(prod[54]),
    .B1(prod[55]),
    .B2(\__uuf__._0818_ ),
    .X(\__uuf__._0415_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0968_ 
  (
    .A(\__uuf__._0817_ ),
    .X(\__uuf__._0343_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0969_ 
  (
    .A(\__uuf__._0811_ ),
    .X(\__uuf__._0819_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0970_ 
  (
    .A(\__uuf__._0813_ ),
    .X(\__uuf__._0820_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0971_ 
  (
    .A1(\__uuf__._0819_ ),
    .A2(\__uuf__._0820_ ),
    .A3(prod[53]),
    .B1(prod[54]),
    .B2(\__uuf__._0818_ ),
    .X(\__uuf__._0414_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0972_ 
  (
    .A(\__uuf__._0817_ ),
    .X(\__uuf__._0342_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0973_ 
  (
    .A1(\__uuf__._0819_ ),
    .A2(\__uuf__._0820_ ),
    .A3(prod[52]),
    .B1(prod[53]),
    .B2(\__uuf__._0818_ ),
    .X(\__uuf__._0413_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0974_ 
  (
    .A(\__uuf__._0817_ ),
    .X(\__uuf__._0341_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0975_ 
  (
    .A1(\__uuf__._0819_ ),
    .A2(\__uuf__._0820_ ),
    .A3(prod[51]),
    .B1(prod[52]),
    .B2(\__uuf__._0818_ ),
    .X(\__uuf__._0412_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0976_ 
  (
    .A(\__uuf__._0817_ ),
    .X(\__uuf__._0340_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0977_ 
  (
    .A1(\__uuf__._0819_ ),
    .A2(\__uuf__._0820_ ),
    .A3(prod[50]),
    .B1(prod[51]),
    .B2(\__uuf__._0818_ ),
    .X(\__uuf__._0411_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0978_ 
  (
    .A(\__uuf__._0816_ ),
    .X(\__uuf__._0821_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0979_ 
  (
    .A(\__uuf__._0821_ ),
    .X(\__uuf__._0339_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0980_ 
  (
    .A(\__uuf__._0774_ ),
    .X(\__uuf__._0822_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0981_ 
  (
    .A1(\__uuf__._0819_ ),
    .A2(\__uuf__._0820_ ),
    .A3(prod[49]),
    .B1(prod[50]),
    .B2(\__uuf__._0822_ ),
    .X(\__uuf__._0410_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0982_ 
  (
    .A(\__uuf__._0821_ ),
    .X(\__uuf__._0338_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0983_ 
  (
    .A(\__uuf__._0811_ ),
    .X(\__uuf__._0823_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0984_ 
  (
    .A(\__uuf__._0813_ ),
    .X(\__uuf__._0824_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0985_ 
  (
    .A1(\__uuf__._0823_ ),
    .A2(\__uuf__._0824_ ),
    .A3(prod[48]),
    .B1(prod[49]),
    .B2(\__uuf__._0822_ ),
    .X(\__uuf__._0409_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0986_ 
  (
    .A(\__uuf__._0821_ ),
    .X(\__uuf__._0337_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0987_ 
  (
    .A1(\__uuf__._0823_ ),
    .A2(\__uuf__._0824_ ),
    .A3(prod[47]),
    .B1(prod[48]),
    .B2(\__uuf__._0822_ ),
    .X(\__uuf__._0408_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0988_ 
  (
    .A(\__uuf__._0821_ ),
    .X(\__uuf__._0336_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0989_ 
  (
    .A1(\__uuf__._0823_ ),
    .A2(\__uuf__._0824_ ),
    .A3(prod[46]),
    .B1(prod[47]),
    .B2(\__uuf__._0822_ ),
    .X(\__uuf__._0407_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0990_ 
  (
    .A(\__uuf__._0821_ ),
    .X(\__uuf__._0335_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0991_ 
  (
    .A1(\__uuf__._0823_ ),
    .A2(\__uuf__._0824_ ),
    .A3(prod[45]),
    .B1(prod[46]),
    .B2(\__uuf__._0822_ ),
    .X(\__uuf__._0406_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0992_ 
  (
    .A(\__uuf__._0816_ ),
    .X(\__uuf__._0825_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0993_ 
  (
    .A(\__uuf__._0825_ ),
    .X(\__uuf__._0334_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0994_ 
  (
    .A(\__uuf__._0773_ ),
    .X(\__uuf__._0826_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0995_ 
  (
    .A(\__uuf__._0826_ ),
    .X(\__uuf__._0827_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._0996_ 
  (
    .A1(\__uuf__._0823_ ),
    .A2(\__uuf__._0824_ ),
    .A3(prod[44]),
    .B1(prod[45]),
    .B2(\__uuf__._0827_ ),
    .X(\__uuf__._0405_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0997_ 
  (
    .A(\__uuf__._0825_ ),
    .X(\__uuf__._0333_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0998_ 
  (
    .A(\__uuf__._0811_ ),
    .X(\__uuf__._0828_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._0999_ 
  (
    .A(\__uuf__._0813_ ),
    .X(\__uuf__._0829_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1000_ 
  (
    .A1(\__uuf__._0828_ ),
    .A2(\__uuf__._0829_ ),
    .A3(prod[43]),
    .B1(prod[44]),
    .B2(\__uuf__._0827_ ),
    .X(\__uuf__._0404_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1001_ 
  (
    .A(\__uuf__._0825_ ),
    .X(\__uuf__._0332_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1002_ 
  (
    .A1(\__uuf__._0828_ ),
    .A2(\__uuf__._0829_ ),
    .A3(prod[42]),
    .B1(prod[43]),
    .B2(\__uuf__._0827_ ),
    .X(\__uuf__._0403_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1003_ 
  (
    .A(\__uuf__._0825_ ),
    .X(\__uuf__._0331_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1004_ 
  (
    .A1(\__uuf__._0828_ ),
    .A2(\__uuf__._0829_ ),
    .A3(prod[41]),
    .B1(prod[42]),
    .B2(\__uuf__._0827_ ),
    .X(\__uuf__._0402_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1005_ 
  (
    .A(\__uuf__._0825_ ),
    .X(\__uuf__._0330_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1006_ 
  (
    .A1(\__uuf__._0828_ ),
    .A2(\__uuf__._0829_ ),
    .A3(prod[40]),
    .B1(prod[41]),
    .B2(\__uuf__._0827_ ),
    .X(\__uuf__._0401_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1007_ 
  (
    .A(\__uuf__._0816_ ),
    .X(\__uuf__._0830_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1008_ 
  (
    .A(\__uuf__._0830_ ),
    .X(\__uuf__._0329_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1009_ 
  (
    .A(\__uuf__._0826_ ),
    .X(\__uuf__._0831_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1010_ 
  (
    .A1(\__uuf__._0828_ ),
    .A2(\__uuf__._0829_ ),
    .A3(prod[39]),
    .B1(prod[40]),
    .B2(\__uuf__._0831_ ),
    .X(\__uuf__._0400_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1011_ 
  (
    .A(\__uuf__._0830_ ),
    .X(\__uuf__._0328_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1012_ 
  (
    .A(\__uuf__._0811_ ),
    .X(\__uuf__._0832_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1013_ 
  (
    .A(\__uuf__._0813_ ),
    .X(\__uuf__._0833_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1014_ 
  (
    .A1(\__uuf__._0832_ ),
    .A2(\__uuf__._0833_ ),
    .A3(prod[38]),
    .B1(prod[39]),
    .B2(\__uuf__._0831_ ),
    .X(\__uuf__._0399_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1015_ 
  (
    .A(\__uuf__._0830_ ),
    .X(\__uuf__._0327_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1016_ 
  (
    .A1(\__uuf__._0832_ ),
    .A2(\__uuf__._0833_ ),
    .A3(prod[37]),
    .B1(prod[38]),
    .B2(\__uuf__._0831_ ),
    .X(\__uuf__._0398_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1017_ 
  (
    .A(\__uuf__._0830_ ),
    .X(\__uuf__._0326_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1018_ 
  (
    .A1(\__uuf__._0832_ ),
    .A2(\__uuf__._0833_ ),
    .A3(prod[36]),
    .B1(prod[37]),
    .B2(\__uuf__._0831_ ),
    .X(\__uuf__._0397_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1019_ 
  (
    .A(\__uuf__._0830_ ),
    .X(\__uuf__._0325_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1020_ 
  (
    .A1(\__uuf__._0832_ ),
    .A2(\__uuf__._0833_ ),
    .A3(prod[35]),
    .B1(prod[36]),
    .B2(\__uuf__._0831_ ),
    .X(\__uuf__._0396_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1021_ 
  (
    .A(\__uuf__._0816_ ),
    .X(\__uuf__._0834_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1022_ 
  (
    .A(\__uuf__._0834_ ),
    .X(\__uuf__._0324_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1023_ 
  (
    .A(\__uuf__._0826_ ),
    .X(\__uuf__._0835_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1024_ 
  (
    .A1(\__uuf__._0832_ ),
    .A2(\__uuf__._0833_ ),
    .A3(prod[34]),
    .B1(prod[35]),
    .B2(\__uuf__._0835_ ),
    .X(\__uuf__._0395_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1025_ 
  (
    .A(\__uuf__._0834_ ),
    .X(\__uuf__._0323_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1026_ 
  (
    .A(\__uuf__._0772_ ),
    .X(\__uuf__._0836_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1027_ 
  (
    .A(\__uuf__._0836_ ),
    .X(\__uuf__._0837_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1028_ 
  (
    .A(\__uuf__._0787_ ),
    .X(\__uuf__._0838_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1029_ 
  (
    .A(\__uuf__._0838_ ),
    .X(\__uuf__._0839_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1030_ 
  (
    .A1(\__uuf__._0837_ ),
    .A2(\__uuf__._0839_ ),
    .A3(prod[33]),
    .B1(prod[34]),
    .B2(\__uuf__._0835_ ),
    .X(\__uuf__._0394_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1031_ 
  (
    .A(\__uuf__._0834_ ),
    .X(\__uuf__._0322_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1032_ 
  (
    .A1(\__uuf__._0837_ ),
    .A2(\__uuf__._0839_ ),
    .A3(prod[32]),
    .B1(prod[33]),
    .B2(\__uuf__._0835_ ),
    .X(\__uuf__._0393_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1033_ 
  (
    .A(\__uuf__._0834_ ),
    .X(\__uuf__._0321_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1034_ 
  (
    .A1(\__uuf__._0837_ ),
    .A2(\__uuf__._0839_ ),
    .A3(prod[31]),
    .B1(prod[32]),
    .B2(\__uuf__._0835_ ),
    .X(\__uuf__._0392_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1035_ 
  (
    .A(\__uuf__._0834_ ),
    .X(\__uuf__._0320_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1036_ 
  (
    .A1(\__uuf__._0837_ ),
    .A2(\__uuf__._0839_ ),
    .A3(prod[30]),
    .B1(prod[31]),
    .B2(\__uuf__._0835_ ),
    .X(\__uuf__._0391_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1037_ 
  (
    .A(\__uuf__._0815_ ),
    .X(\__uuf__._0840_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1038_ 
  (
    .A(\__uuf__._0840_ ),
    .X(\__uuf__._0841_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1039_ 
  (
    .A(\__uuf__._0841_ ),
    .X(\__uuf__._0319_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1040_ 
  (
    .A(\__uuf__._0826_ ),
    .X(\__uuf__._0842_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1041_ 
  (
    .A1(\__uuf__._0837_ ),
    .A2(\__uuf__._0839_ ),
    .A3(prod[29]),
    .B1(prod[30]),
    .B2(\__uuf__._0842_ ),
    .X(\__uuf__._0390_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1042_ 
  (
    .A(\__uuf__._0841_ ),
    .X(\__uuf__._0318_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1043_ 
  (
    .A(\__uuf__._0836_ ),
    .X(\__uuf__._0843_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1044_ 
  (
    .A(\__uuf__._0838_ ),
    .X(\__uuf__._0844_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1045_ 
  (
    .A1(\__uuf__._0843_ ),
    .A2(\__uuf__._0844_ ),
    .A3(prod[28]),
    .B1(prod[29]),
    .B2(\__uuf__._0842_ ),
    .X(\__uuf__._0389_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1046_ 
  (
    .A(\__uuf__._0841_ ),
    .X(\__uuf__._0317_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1047_ 
  (
    .A1(\__uuf__._0843_ ),
    .A2(\__uuf__._0844_ ),
    .A3(prod[27]),
    .B1(prod[28]),
    .B2(\__uuf__._0842_ ),
    .X(\__uuf__._0388_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1048_ 
  (
    .A(\__uuf__._0841_ ),
    .X(\__uuf__._0316_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1049_ 
  (
    .A1(\__uuf__._0843_ ),
    .A2(\__uuf__._0844_ ),
    .A3(prod[26]),
    .B1(prod[27]),
    .B2(\__uuf__._0842_ ),
    .X(\__uuf__._0387_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1050_ 
  (
    .A(\__uuf__._0841_ ),
    .X(\__uuf__._0315_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1051_ 
  (
    .A1(\__uuf__._0843_ ),
    .A2(\__uuf__._0844_ ),
    .A3(prod[25]),
    .B1(prod[26]),
    .B2(\__uuf__._0842_ ),
    .X(\__uuf__._0386_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1052_ 
  (
    .A(\__uuf__._0840_ ),
    .X(\__uuf__._0845_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1053_ 
  (
    .A(\__uuf__._0845_ ),
    .X(\__uuf__._0314_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1054_ 
  (
    .A(\__uuf__._0826_ ),
    .X(\__uuf__._0846_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1055_ 
  (
    .A1(\__uuf__._0843_ ),
    .A2(\__uuf__._0844_ ),
    .A3(prod[24]),
    .B1(prod[25]),
    .B2(\__uuf__._0846_ ),
    .X(\__uuf__._0385_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1056_ 
  (
    .A(\__uuf__._0845_ ),
    .X(\__uuf__._0313_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1057_ 
  (
    .A(\__uuf__._0836_ ),
    .X(\__uuf__._0847_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1058_ 
  (
    .A(\__uuf__._0838_ ),
    .X(\__uuf__._0848_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1059_ 
  (
    .A1(\__uuf__._0847_ ),
    .A2(\__uuf__._0848_ ),
    .A3(prod[23]),
    .B1(prod[24]),
    .B2(\__uuf__._0846_ ),
    .X(\__uuf__._0384_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1060_ 
  (
    .A(\__uuf__._0845_ ),
    .X(\__uuf__._0312_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1061_ 
  (
    .A1(\__uuf__._0847_ ),
    .A2(\__uuf__._0848_ ),
    .A3(prod[22]),
    .B1(prod[23]),
    .B2(\__uuf__._0846_ ),
    .X(\__uuf__._0383_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1062_ 
  (
    .A(\__uuf__._0845_ ),
    .X(\__uuf__._0311_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1063_ 
  (
    .A1(\__uuf__._0847_ ),
    .A2(\__uuf__._0848_ ),
    .A3(prod[21]),
    .B1(prod[22]),
    .B2(\__uuf__._0846_ ),
    .X(\__uuf__._0382_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1064_ 
  (
    .A(\__uuf__._0845_ ),
    .X(\__uuf__._0310_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1065_ 
  (
    .A1(\__uuf__._0847_ ),
    .A2(\__uuf__._0848_ ),
    .A3(prod[20]),
    .B1(prod[21]),
    .B2(\__uuf__._0846_ ),
    .X(\__uuf__._0381_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1066_ 
  (
    .A(\__uuf__._0840_ ),
    .X(\__uuf__._0849_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1067_ 
  (
    .A(\__uuf__._0849_ ),
    .X(\__uuf__._0309_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1068_ 
  (
    .A(\__uuf__._0803_ ),
    .X(\__uuf__._0850_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1069_ 
  (
    .A1(\__uuf__._0847_ ),
    .A2(\__uuf__._0848_ ),
    .A3(prod[19]),
    .B1(prod[20]),
    .B2(\__uuf__._0850_ ),
    .X(\__uuf__._0380_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1070_ 
  (
    .A(\__uuf__._0849_ ),
    .X(\__uuf__._0308_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1071_ 
  (
    .A(\__uuf__._0836_ ),
    .X(\__uuf__._0851_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1072_ 
  (
    .A(\__uuf__._0838_ ),
    .X(\__uuf__._0852_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1073_ 
  (
    .A1(\__uuf__._0851_ ),
    .A2(\__uuf__._0852_ ),
    .A3(prod[18]),
    .B1(prod[19]),
    .B2(\__uuf__._0850_ ),
    .X(\__uuf__._0379_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1074_ 
  (
    .A(\__uuf__._0849_ ),
    .X(\__uuf__._0307_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1075_ 
  (
    .A1(\__uuf__._0851_ ),
    .A2(\__uuf__._0852_ ),
    .A3(prod[17]),
    .B1(prod[18]),
    .B2(\__uuf__._0850_ ),
    .X(\__uuf__._0378_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1076_ 
  (
    .A(\__uuf__._0849_ ),
    .X(\__uuf__._0306_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1077_ 
  (
    .A1(\__uuf__._0851_ ),
    .A2(\__uuf__._0852_ ),
    .A3(prod[16]),
    .B1(prod[17]),
    .B2(\__uuf__._0850_ ),
    .X(\__uuf__._0377_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1078_ 
  (
    .A(\__uuf__._0849_ ),
    .X(\__uuf__._0305_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1079_ 
  (
    .A1(\__uuf__._0851_ ),
    .A2(\__uuf__._0852_ ),
    .A3(prod[15]),
    .B1(prod[16]),
    .B2(\__uuf__._0850_ ),
    .X(\__uuf__._0376_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1080_ 
  (
    .A(\__uuf__._0840_ ),
    .X(\__uuf__._0853_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1081_ 
  (
    .A(\__uuf__._0853_ ),
    .X(\__uuf__._0304_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1082_ 
  (
    .A(\__uuf__._0803_ ),
    .X(\__uuf__._0854_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1083_ 
  (
    .A1(\__uuf__._0851_ ),
    .A2(\__uuf__._0852_ ),
    .A3(prod[14]),
    .B1(prod[15]),
    .B2(\__uuf__._0854_ ),
    .X(\__uuf__._0375_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1084_ 
  (
    .A(\__uuf__._0853_ ),
    .X(\__uuf__._0303_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1085_ 
  (
    .A(\__uuf__._0836_ ),
    .X(\__uuf__._0855_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1086_ 
  (
    .A(\__uuf__._0838_ ),
    .X(\__uuf__._0856_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1087_ 
  (
    .A1(\__uuf__._0855_ ),
    .A2(\__uuf__._0856_ ),
    .A3(prod[13]),
    .B1(prod[14]),
    .B2(\__uuf__._0854_ ),
    .X(\__uuf__._0374_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1088_ 
  (
    .A(\__uuf__._0853_ ),
    .X(\__uuf__._0302_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1089_ 
  (
    .A1(\__uuf__._0855_ ),
    .A2(\__uuf__._0856_ ),
    .A3(prod[12]),
    .B1(prod[13]),
    .B2(\__uuf__._0854_ ),
    .X(\__uuf__._0373_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1090_ 
  (
    .A(\__uuf__._0853_ ),
    .X(\__uuf__._0301_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1091_ 
  (
    .A1(\__uuf__._0855_ ),
    .A2(\__uuf__._0856_ ),
    .A3(prod[11]),
    .B1(prod[12]),
    .B2(\__uuf__._0854_ ),
    .X(\__uuf__._0372_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1092_ 
  (
    .A(\__uuf__._0853_ ),
    .X(\__uuf__._0300_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1093_ 
  (
    .A1(\__uuf__._0855_ ),
    .A2(\__uuf__._0856_ ),
    .A3(prod[10]),
    .B1(prod[11]),
    .B2(\__uuf__._0854_ ),
    .X(\__uuf__._0371_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1094_ 
  (
    .A(\__uuf__._0840_ ),
    .X(\__uuf__._0857_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1095_ 
  (
    .A(\__uuf__._0857_ ),
    .X(\__uuf__._0299_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1096_ 
  (
    .A(\__uuf__._0803_ ),
    .X(\__uuf__._0858_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1097_ 
  (
    .A1(\__uuf__._0855_ ),
    .A2(\__uuf__._0856_ ),
    .A3(prod[9]),
    .B1(prod[10]),
    .B2(\__uuf__._0858_ ),
    .X(\__uuf__._0370_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1098_ 
  (
    .A(\__uuf__._0857_ ),
    .X(\__uuf__._0298_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1099_ 
  (
    .A(\__uuf__._0772_ ),
    .X(\__uuf__._0859_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1100_ 
  (
    .A(\__uuf__._0787_ ),
    .X(\__uuf__._0860_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1101_ 
  (
    .A(\__uuf__._0860_ ),
    .X(\__uuf__._0861_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1102_ 
  (
    .A1(\__uuf__._0859_ ),
    .A2(\__uuf__._0861_ ),
    .A3(prod[8]),
    .B1(prod[9]),
    .B2(\__uuf__._0858_ ),
    .X(\__uuf__._0369_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1103_ 
  (
    .A(\__uuf__._0857_ ),
    .X(\__uuf__._0297_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1104_ 
  (
    .A1(\__uuf__._0859_ ),
    .A2(\__uuf__._0861_ ),
    .A3(prod[7]),
    .B1(prod[8]),
    .B2(\__uuf__._0858_ ),
    .X(\__uuf__._0368_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1105_ 
  (
    .A(\__uuf__._0857_ ),
    .X(\__uuf__._0296_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1106_ 
  (
    .A1(\__uuf__._0859_ ),
    .A2(\__uuf__._0861_ ),
    .A3(prod[6]),
    .B1(prod[7]),
    .B2(\__uuf__._0858_ ),
    .X(\__uuf__._0367_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1107_ 
  (
    .A(\__uuf__._0857_ ),
    .X(\__uuf__._0295_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1108_ 
  (
    .A1(\__uuf__._0859_ ),
    .A2(\__uuf__._0861_ ),
    .A3(prod[5]),
    .B1(prod[6]),
    .B2(\__uuf__._0858_ ),
    .X(\__uuf__._0366_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1109_ 
  (
    .A(\__uuf__._0815_ ),
    .X(\__uuf__._0862_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1110_ 
  (
    .A(\__uuf__._0862_ ),
    .X(\__uuf__._0863_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1111_ 
  (
    .A(\__uuf__._0863_ ),
    .X(\__uuf__._0294_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1112_ 
  (
    .A(\__uuf__._0803_ ),
    .X(\__uuf__._0864_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1113_ 
  (
    .A1(\__uuf__._0859_ ),
    .A2(\__uuf__._0861_ ),
    .A3(prod[4]),
    .B1(prod[5]),
    .B2(\__uuf__._0864_ ),
    .X(\__uuf__._0365_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1114_ 
  (
    .A(\__uuf__._0863_ ),
    .X(\__uuf__._0293_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1115_ 
  (
    .A(\__uuf__._0860_ ),
    .X(\__uuf__._0865_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1116_ 
  (
    .A1(\__uuf__._0805_ ),
    .A2(\__uuf__._0865_ ),
    .A3(prod[3]),
    .B1(prod[4]),
    .B2(\__uuf__._0864_ ),
    .X(\__uuf__._0364_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1117_ 
  (
    .A(\__uuf__._0863_ ),
    .X(\__uuf__._0292_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1118_ 
  (
    .A1(\__uuf__._0805_ ),
    .A2(\__uuf__._0865_ ),
    .A3(prod[2]),
    .B1(prod[3]),
    .B2(\__uuf__._0864_ ),
    .X(\__uuf__._0363_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1119_ 
  (
    .A(\__uuf__._0863_ ),
    .X(\__uuf__._0291_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1120_ 
  (
    .A1(\__uuf__._0805_ ),
    .A2(\__uuf__._0865_ ),
    .A3(prod[1]),
    .B1(prod[2]),
    .B2(\__uuf__._0864_ ),
    .X(\__uuf__._0362_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1121_ 
  (
    .A(\__uuf__._0863_ ),
    .X(\__uuf__._0290_ )
  );


  sky130_fd_sc_hd__a32o_4
  \__uuf__._1122_ 
  (
    .A1(\__uuf__._0805_ ),
    .A2(\__uuf__._0865_ ),
    .A3(prod[0]),
    .B1(prod[1]),
    .B2(\__uuf__._0864_ ),
    .X(\__uuf__._0361_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1123_ 
  (
    .A(\__uuf__._0862_ ),
    .X(\__uuf__._0866_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1124_ 
  (
    .A(\__uuf__._0866_ ),
    .X(\__uuf__._0289_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1125_ 
  (
    .A(\__uuf__._0866_ ),
    .X(\__uuf__._0288_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1126_ 
  (
    .A(\__uuf__._0866_ ),
    .X(\__uuf__._0287_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1127_ 
  (
    .A(\__uuf__._0866_ ),
    .X(\__uuf__._0286_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1128_ 
  (
    .A(\__uuf__._0866_ ),
    .X(\__uuf__._0285_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1129_ 
  (
    .A(\__uuf__._0862_ ),
    .X(\__uuf__._0867_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1130_ 
  (
    .A(\__uuf__._0867_ ),
    .X(\__uuf__._0284_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1131_ 
  (
    .A(\__uuf__._0867_ ),
    .X(\__uuf__._0283_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1132_ 
  (
    .A(\__uuf__._0867_ ),
    .X(\__uuf__._0282_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1133_ 
  (
    .A(\__uuf__._0867_ ),
    .X(\__uuf__._0281_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1134_ 
  (
    .A(\__uuf__._0867_ ),
    .X(\__uuf__._0280_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1135_ 
  (
    .A(\__uuf__._0862_ ),
    .X(\__uuf__._0868_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1136_ 
  (
    .A(\__uuf__._0868_ ),
    .X(\__uuf__._0279_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1137_ 
  (
    .A(\__uuf__._0868_ ),
    .X(\__uuf__._0278_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1138_ 
  (
    .A(\__uuf__._0868_ ),
    .X(\__uuf__._0277_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1139_ 
  (
    .A(\__uuf__._0868_ ),
    .X(\__uuf__._0276_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1140_ 
  (
    .A(\__uuf__._0868_ ),
    .X(\__uuf__._0275_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1141_ 
  (
    .A(\__uuf__._0862_ ),
    .X(\__uuf__._0869_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1142_ 
  (
    .A(\__uuf__._0869_ ),
    .X(\__uuf__._0274_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1143_ 
  (
    .A(\__uuf__._0869_ ),
    .X(\__uuf__._0273_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1144_ 
  (
    .A(\__uuf__._0869_ ),
    .X(\__uuf__._0272_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1145_ 
  (
    .A(\__uuf__._0869_ ),
    .X(\__uuf__._0271_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1146_ 
  (
    .A(\__uuf__._0869_ ),
    .X(\__uuf__._0270_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1147_ 
  (
    .A(\__uuf__._0793_ ),
    .X(\__uuf__._0870_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1148_ 
  (
    .A(\__uuf__._0870_ ),
    .X(\__uuf__._0871_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1149_ 
  (
    .A(\__uuf__._0871_ ),
    .X(\__uuf__._0269_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1150_ 
  (
    .A(\__uuf__._0871_ ),
    .X(\__uuf__._0268_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1151_ 
  (
    .A(\__uuf__._0871_ ),
    .X(\__uuf__._0267_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1152_ 
  (
    .A(\__uuf__._0871_ ),
    .X(\__uuf__._0266_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1153_ 
  (
    .A(\__uuf__._0871_ ),
    .X(\__uuf__._0265_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1154_ 
  (
    .A(\__uuf__._0870_ ),
    .X(\__uuf__._0872_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1155_ 
  (
    .A(\__uuf__._0872_ ),
    .X(\__uuf__._0264_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1156_ 
  (
    .A(\__uuf__._0872_ ),
    .X(\__uuf__._0263_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1157_ 
  (
    .A(\__uuf__._0872_ ),
    .X(\__uuf__._0262_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1158_ 
  (
    .A(\__uuf__._0872_ ),
    .X(\__uuf__._0261_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1159_ 
  (
    .A(\__uuf__._0872_ ),
    .X(\__uuf__._0260_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1160_ 
  (
    .A(\__uuf__._0870_ ),
    .X(\__uuf__._0873_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1161_ 
  (
    .A(\__uuf__._0873_ ),
    .X(\__uuf__._0259_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1162_ 
  (
    .A(\__uuf__._0873_ ),
    .X(\__uuf__._0258_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1163_ 
  (
    .A(\__uuf__._0873_ ),
    .X(\__uuf__._0257_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1164_ 
  (
    .A(\__uuf__._0873_ ),
    .X(\__uuf__._0256_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1165_ 
  (
    .A(\__uuf__._0873_ ),
    .X(\__uuf__._0255_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1166_ 
  (
    .A(\__uuf__._0870_ ),
    .X(\__uuf__._0874_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1167_ 
  (
    .A(\__uuf__._0874_ ),
    .X(\__uuf__._0254_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1168_ 
  (
    .A(\__uuf__._0874_ ),
    .X(\__uuf__._0253_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1169_ 
  (
    .A(\__uuf__._0874_ ),
    .X(\__uuf__._0252_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1170_ 
  (
    .A(\__uuf__._0874_ ),
    .X(\__uuf__._0251_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1171_ 
  (
    .A(\__uuf__._0874_ ),
    .X(\__uuf__._0250_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1172_ 
  (
    .A(\__uuf__._0870_ ),
    .X(\__uuf__._0875_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1173_ 
  (
    .A(\__uuf__._0875_ ),
    .X(\__uuf__._0249_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1174_ 
  (
    .A(\__uuf__._0875_ ),
    .X(\__uuf__._0248_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1175_ 
  (
    .A(\__uuf__._0875_ ),
    .X(\__uuf__._0247_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1176_ 
  (
    .A(\__uuf__._0875_ ),
    .X(\__uuf__._0246_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1177_ 
  (
    .A(\__uuf__._0875_ ),
    .X(\__uuf__._0245_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1178_ 
  (
    .A(\__uuf__._0793_ ),
    .X(\__uuf__._0876_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1179_ 
  (
    .A(\__uuf__._0876_ ),
    .X(\__uuf__._0877_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1180_ 
  (
    .A(\__uuf__._0877_ ),
    .X(\__uuf__._0244_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1181_ 
  (
    .A(\__uuf__._0877_ ),
    .X(\__uuf__._0243_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1182_ 
  (
    .A(\__uuf__._0877_ ),
    .X(\__uuf__._0242_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1183_ 
  (
    .A(\__uuf__._0877_ ),
    .X(\__uuf__._0241_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1184_ 
  (
    .A(\__uuf__._0877_ ),
    .X(\__uuf__._0240_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1185_ 
  (
    .A(\__uuf__._0876_ ),
    .X(\__uuf__._0878_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1186_ 
  (
    .A(\__uuf__._0878_ ),
    .X(\__uuf__._0239_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1187_ 
  (
    .A(\__uuf__._0878_ ),
    .X(\__uuf__._0238_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1188_ 
  (
    .A(\__uuf__._0878_ ),
    .X(\__uuf__._0237_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1189_ 
  (
    .A(\__uuf__._0878_ ),
    .X(\__uuf__._0236_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1190_ 
  (
    .A(\__uuf__._0878_ ),
    .X(\__uuf__._0235_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1191_ 
  (
    .A(\__uuf__._0876_ ),
    .X(\__uuf__._0879_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1192_ 
  (
    .A(\__uuf__._0879_ ),
    .X(\__uuf__._0234_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1193_ 
  (
    .A(\__uuf__._0879_ ),
    .X(\__uuf__._0233_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1194_ 
  (
    .A(\__uuf__._0879_ ),
    .X(\__uuf__._0232_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1195_ 
  (
    .A(\__uuf__._0879_ ),
    .X(\__uuf__._0231_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1196_ 
  (
    .A(\__uuf__._0879_ ),
    .X(\__uuf__._0230_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1197_ 
  (
    .A(\__uuf__._0876_ ),
    .X(\__uuf__._0880_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1198_ 
  (
    .A(\__uuf__._0880_ ),
    .X(\__uuf__._0229_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1199_ 
  (
    .A(\__uuf__._0880_ ),
    .X(\__uuf__._0228_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1200_ 
  (
    .A(\__uuf__._0880_ ),
    .X(\__uuf__._0227_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1201_ 
  (
    .A(\__uuf__._0880_ ),
    .X(\__uuf__._0226_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1202_ 
  (
    .A(\__uuf__._0880_ ),
    .X(\__uuf__._0225_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1203_ 
  (
    .A(\__uuf__._0876_ ),
    .X(\__uuf__._0881_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1204_ 
  (
    .A(\__uuf__._0881_ ),
    .X(\__uuf__._0224_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1205_ 
  (
    .A(\__uuf__._0881_ ),
    .X(\__uuf__._0223_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1206_ 
  (
    .A(\__uuf__._0881_ ),
    .X(\__uuf__._0222_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1207_ 
  (
    .A(\__uuf__._0881_ ),
    .X(\__uuf__._0221_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1208_ 
  (
    .A(\__uuf__._0881_ ),
    .X(\__uuf__._0220_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1209_ 
  (
    .A(\__uuf__._0793_ ),
    .X(\__uuf__._0432_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1210_ 
  (
    .A(\__uuf__._0432_ ),
    .X(\__uuf__._0433_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1211_ 
  (
    .A(\__uuf__._0433_ ),
    .X(\__uuf__._0219_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1212_ 
  (
    .A(\__uuf__._0433_ ),
    .X(\__uuf__._0218_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1213_ 
  (
    .A(\__uuf__._0433_ ),
    .X(\__uuf__._0217_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1214_ 
  (
    .A(\__uuf__._0433_ ),
    .X(\__uuf__._0216_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1215_ 
  (
    .A(\__uuf__._0433_ ),
    .X(\__uuf__._0215_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1216_ 
  (
    .A(\__uuf__._0432_ ),
    .X(\__uuf__._0434_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1217_ 
  (
    .A(\__uuf__._0434_ ),
    .X(\__uuf__._0214_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1218_ 
  (
    .A(\__uuf__._0434_ ),
    .X(\__uuf__._0213_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1219_ 
  (
    .A(\__uuf__._0434_ ),
    .X(\__uuf__._0212_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1220_ 
  (
    .A(\__uuf__._0434_ ),
    .X(\__uuf__._0211_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1221_ 
  (
    .A(\__uuf__._0434_ ),
    .X(\__uuf__._0210_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1222_ 
  (
    .A(\__uuf__._0432_ ),
    .X(\__uuf__._0435_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1223_ 
  (
    .A(\__uuf__._0435_ ),
    .X(\__uuf__._0209_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1224_ 
  (
    .A(\__uuf__._0435_ ),
    .X(\__uuf__._0208_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1225_ 
  (
    .A(\__uuf__._0435_ ),
    .X(\__uuf__._0207_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1226_ 
  (
    .A(\__uuf__._0435_ ),
    .X(\__uuf__._0206_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1227_ 
  (
    .A(\__uuf__._0435_ ),
    .X(\__uuf__._0205_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1228_ 
  (
    .A(\__uuf__._0432_ ),
    .X(\__uuf__._0436_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1229_ 
  (
    .A(\__uuf__._0436_ ),
    .X(\__uuf__._0204_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1230_ 
  (
    .A(\__uuf__._0436_ ),
    .X(\__uuf__._0203_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1231_ 
  (
    .A(\__uuf__._0436_ ),
    .X(\__uuf__._0202_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1232_ 
  (
    .A(\__uuf__._0436_ ),
    .X(\__uuf__._0201_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1233_ 
  (
    .A(\__uuf__._0436_ ),
    .X(\__uuf__._0200_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1234_ 
  (
    .A(\__uuf__._0432_ ),
    .X(\__uuf__._0437_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1235_ 
  (
    .A(\__uuf__._0437_ ),
    .X(\__uuf__._0199_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1236_ 
  (
    .A(\__uuf__._0437_ ),
    .X(\__uuf__._0198_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1237_ 
  (
    .A(\__uuf__._0437_ ),
    .X(\__uuf__._0197_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1238_ 
  (
    .A(\__uuf__._0437_ ),
    .X(\__uuf__._0196_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1239_ 
  (
    .A(\__uuf__._0437_ ),
    .X(\__uuf__._0195_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1240_ 
  (
    .A(\__uuf__._0793_ ),
    .X(\__uuf__._0438_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1241_ 
  (
    .A(\__uuf__._0438_ ),
    .X(\__uuf__._0439_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1242_ 
  (
    .A(\__uuf__._0439_ ),
    .X(\__uuf__._0194_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1243_ 
  (
    .A(\__uuf__._0439_ ),
    .X(\__uuf__._0193_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1244_ 
  (
    .A(\__uuf__._0439_ ),
    .X(\__uuf__._0192_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1245_ 
  (
    .A(\__uuf__._0439_ ),
    .X(\__uuf__._0191_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1246_ 
  (
    .A(\__uuf__._0439_ ),
    .X(\__uuf__._0190_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1247_ 
  (
    .A(\__uuf__._0438_ ),
    .X(\__uuf__._0440_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1248_ 
  (
    .A(\__uuf__._0440_ ),
    .X(\__uuf__._0189_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1249_ 
  (
    .A(\__uuf__._0440_ ),
    .X(\__uuf__._0188_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1250_ 
  (
    .A(\__uuf__._0440_ ),
    .X(\__uuf__._0187_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1251_ 
  (
    .A(\__uuf__._0440_ ),
    .X(\__uuf__._0186_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1252_ 
  (
    .A(\__uuf__._0440_ ),
    .X(\__uuf__._0185_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1253_ 
  (
    .A(\__uuf__._0438_ ),
    .X(\__uuf__._0441_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1254_ 
  (
    .A(\__uuf__._0441_ ),
    .X(\__uuf__._0184_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1255_ 
  (
    .A(\__uuf__._0441_ ),
    .X(\__uuf__._0183_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1256_ 
  (
    .A(\__uuf__._0441_ ),
    .X(\__uuf__._0182_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1257_ 
  (
    .A(\__uuf__._0441_ ),
    .X(\__uuf__._0181_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1258_ 
  (
    .A(\__uuf__._0441_ ),
    .X(\__uuf__._0180_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1259_ 
  (
    .A(\__uuf__._0438_ ),
    .X(\__uuf__._0442_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1260_ 
  (
    .A(\__uuf__._0442_ ),
    .X(\__uuf__._0179_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1261_ 
  (
    .A(\__uuf__._0442_ ),
    .X(\__uuf__._0178_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1262_ 
  (
    .A(\__uuf__._0442_ ),
    .X(\__uuf__._0177_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1263_ 
  (
    .A(\__uuf__._0442_ ),
    .X(\__uuf__._0176_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1264_ 
  (
    .A(\__uuf__._0442_ ),
    .X(\__uuf__._0175_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1265_ 
  (
    .A(\__uuf__._0438_ ),
    .X(\__uuf__._0443_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1266_ 
  (
    .A(\__uuf__._0443_ ),
    .X(\__uuf__._0174_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1267_ 
  (
    .A(\__uuf__._0443_ ),
    .X(\__uuf__._0173_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1268_ 
  (
    .A(\__uuf__._0443_ ),
    .X(\__uuf__._0172_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1269_ 
  (
    .A(\__uuf__._0443_ ),
    .X(\__uuf__._0171_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1270_ 
  (
    .A(\__uuf__._0443_ ),
    .X(\__uuf__._0170_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1271_ 
  (
    .A(\__uuf__._0815_ ),
    .X(\__uuf__._0444_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1272_ 
  (
    .A(\__uuf__._0444_ ),
    .X(\__uuf__._0169_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1273_ 
  (
    .A(\__uuf__._0444_ ),
    .X(\__uuf__._0168_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1274_ 
  (
    .A(\__uuf__._0444_ ),
    .X(\__uuf__._0167_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1275_ 
  (
    .A(\__uuf__._0444_ ),
    .X(\__uuf__._0166_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1276_ 
  (
    .A(\__uuf__._0444_ ),
    .X(\__uuf__._0165_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1277_ 
  (
    .A(\__uuf__._0815_ ),
    .X(\__uuf__._0445_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1278_ 
  (
    .A(\__uuf__._0445_ ),
    .X(\__uuf__._0164_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1279_ 
  (
    .A(\__uuf__._0445_ ),
    .X(\__uuf__._0163_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1280_ 
  (
    .A(\__uuf__._0445_ ),
    .X(\__uuf__._0162_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1281_ 
  (
    .A(\__uuf__._0445_ ),
    .X(\__uuf__._0161_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1282_ 
  (
    .A(\__uuf__._0445_ ),
    .X(\__uuf__._0160_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1283_ 
  (
    .A(\__uuf__._0794_ ),
    .X(\__uuf__._0159_ )
  );


  sky130_fd_sc_hd__and2_4
  \__uuf__._1284_ 
  (
    .A(\__uuf__._0766_ ),
    .B(\__uuf__.fsm.state[1] ),
    .X(\__uuf__._0446_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1285_ 
  (
    .A(\__uuf__._0446_ ),
    .X(done)
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1286_ 
  (
    .A(\__uuf__._0807_ ),
    .X(\__uuf__._0447_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1287_ 
  (
    .A(\__uuf__._0788_ ),
    .X(\__uuf__._0448_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1288_ 
  (
    .A(\__uuf__._0448_ ),
    .X(\__uuf__._0449_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1289_ 
  (
    .A(\__uuf__._0449_ ),
    .X(\__uuf__._0450_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1290_ 
  (
    .A1(\__BoundaryScanRegister_input_32__.dout ),
    .A2(\__uuf__._0447_ ),
    .B1(\__uuf__.shifter.shiftreg[1] ),
    .B2(\__uuf__._0450_ ),
    .X(\__uuf__._0095_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1291_ 
  (
    .A1(\__BoundaryScanRegister_input_33__.dout ),
    .A2(\__uuf__._0447_ ),
    .B1(\__uuf__.shifter.shiftreg[2] ),
    .B2(\__uuf__._0450_ ),
    .X(\__uuf__._0106_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1292_ 
  (
    .A(\__uuf__._0860_ ),
    .X(\__uuf__._0451_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1293_ 
  (
    .A(\__uuf__._0451_ ),
    .X(\__uuf__._0452_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1294_ 
  (
    .A1(\__BoundaryScanRegister_input_34__.dout ),
    .A2(\__uuf__._0452_ ),
    .B1(\__uuf__.shifter.shiftreg[3] ),
    .B2(\__uuf__._0450_ ),
    .X(\__uuf__._0117_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1295_ 
  (
    .A1(\__BoundaryScanRegister_input_35__.dout ),
    .A2(\__uuf__._0452_ ),
    .B1(\__uuf__.shifter.shiftreg[4] ),
    .B2(\__uuf__._0450_ ),
    .X(\__uuf__._0128_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1296_ 
  (
    .A1(\__BoundaryScanRegister_input_36__.dout ),
    .A2(\__uuf__._0452_ ),
    .B1(\__uuf__.shifter.shiftreg[5] ),
    .B2(\__uuf__._0450_ ),
    .X(\__uuf__._0139_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1297_ 
  (
    .A(\__uuf__._0449_ ),
    .X(\__uuf__._0453_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1298_ 
  (
    .A1(\__BoundaryScanRegister_input_37__.dout ),
    .A2(\__uuf__._0452_ ),
    .B1(\__uuf__.shifter.shiftreg[6] ),
    .B2(\__uuf__._0453_ ),
    .X(\__uuf__._0150_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1299_ 
  (
    .A1(\__BoundaryScanRegister_input_38__.dout ),
    .A2(\__uuf__._0452_ ),
    .B1(\__uuf__.shifter.shiftreg[7] ),
    .B2(\__uuf__._0453_ ),
    .X(\__uuf__._0155_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1300_ 
  (
    .A(\__uuf__._0451_ ),
    .X(\__uuf__._0454_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1301_ 
  (
    .A1(\__BoundaryScanRegister_input_39__.dout ),
    .A2(\__uuf__._0454_ ),
    .B1(\__uuf__.shifter.shiftreg[8] ),
    .B2(\__uuf__._0453_ ),
    .X(\__uuf__._0156_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1302_ 
  (
    .A1(\__BoundaryScanRegister_input_40__.dout ),
    .A2(\__uuf__._0454_ ),
    .B1(\__uuf__.shifter.shiftreg[9] ),
    .B2(\__uuf__._0453_ ),
    .X(\__uuf__._0157_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1303_ 
  (
    .A1(\__BoundaryScanRegister_input_41__.dout ),
    .A2(\__uuf__._0454_ ),
    .B1(\__uuf__.shifter.shiftreg[10] ),
    .B2(\__uuf__._0453_ ),
    .X(\__uuf__._0158_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1304_ 
  (
    .A(\__uuf__._0449_ ),
    .X(\__uuf__._0455_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1305_ 
  (
    .A1(\__BoundaryScanRegister_input_42__.dout ),
    .A2(\__uuf__._0454_ ),
    .B1(\__uuf__.shifter.shiftreg[11] ),
    .B2(\__uuf__._0455_ ),
    .X(\__uuf__._0096_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1306_ 
  (
    .A1(\__BoundaryScanRegister_input_43__.dout ),
    .A2(\__uuf__._0454_ ),
    .B1(\__uuf__.shifter.shiftreg[12] ),
    .B2(\__uuf__._0455_ ),
    .X(\__uuf__._0097_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1307_ 
  (
    .A(\__uuf__._0451_ ),
    .X(\__uuf__._0456_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1308_ 
  (
    .A1(\__BoundaryScanRegister_input_44__.dout ),
    .A2(\__uuf__._0456_ ),
    .B1(\__uuf__.shifter.shiftreg[13] ),
    .B2(\__uuf__._0455_ ),
    .X(\__uuf__._0098_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1309_ 
  (
    .A1(\__BoundaryScanRegister_input_45__.dout ),
    .A2(\__uuf__._0456_ ),
    .B1(\__uuf__.shifter.shiftreg[14] ),
    .B2(\__uuf__._0455_ ),
    .X(\__uuf__._0099_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1310_ 
  (
    .A1(\__BoundaryScanRegister_input_46__.dout ),
    .A2(\__uuf__._0456_ ),
    .B1(\__uuf__.shifter.shiftreg[15] ),
    .B2(\__uuf__._0455_ ),
    .X(\__uuf__._0100_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1311_ 
  (
    .A(\__uuf__._0788_ ),
    .X(\__uuf__._0457_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1312_ 
  (
    .A(\__uuf__._0457_ ),
    .X(\__uuf__._0458_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1313_ 
  (
    .A1(\__BoundaryScanRegister_input_47__.dout ),
    .A2(\__uuf__._0456_ ),
    .B1(\__uuf__.shifter.shiftreg[16] ),
    .B2(\__uuf__._0458_ ),
    .X(\__uuf__._0101_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1314_ 
  (
    .A1(\__BoundaryScanRegister_input_48__.dout ),
    .A2(\__uuf__._0456_ ),
    .B1(\__uuf__.shifter.shiftreg[17] ),
    .B2(\__uuf__._0458_ ),
    .X(\__uuf__._0102_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1315_ 
  (
    .A(\__uuf__._0451_ ),
    .X(\__uuf__._0459_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1316_ 
  (
    .A1(\__BoundaryScanRegister_input_49__.dout ),
    .A2(\__uuf__._0459_ ),
    .B1(\__uuf__.shifter.shiftreg[18] ),
    .B2(\__uuf__._0458_ ),
    .X(\__uuf__._0103_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1317_ 
  (
    .A1(\__BoundaryScanRegister_input_50__.dout ),
    .A2(\__uuf__._0459_ ),
    .B1(\__uuf__.shifter.shiftreg[19] ),
    .B2(\__uuf__._0458_ ),
    .X(\__uuf__._0104_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1318_ 
  (
    .A1(\__BoundaryScanRegister_input_51__.dout ),
    .A2(\__uuf__._0459_ ),
    .B1(\__uuf__.shifter.shiftreg[20] ),
    .B2(\__uuf__._0458_ ),
    .X(\__uuf__._0105_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1319_ 
  (
    .A(\__uuf__._0457_ ),
    .X(\__uuf__._0460_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1320_ 
  (
    .A1(\__BoundaryScanRegister_input_52__.dout ),
    .A2(\__uuf__._0459_ ),
    .B1(\__uuf__.shifter.shiftreg[21] ),
    .B2(\__uuf__._0460_ ),
    .X(\__uuf__._0107_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1321_ 
  (
    .A1(\__BoundaryScanRegister_input_53__.dout ),
    .A2(\__uuf__._0459_ ),
    .B1(\__uuf__.shifter.shiftreg[22] ),
    .B2(\__uuf__._0460_ ),
    .X(\__uuf__._0108_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1322_ 
  (
    .A(\__uuf__._0451_ ),
    .X(\__uuf__._0461_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1323_ 
  (
    .A1(\__BoundaryScanRegister_input_54__.dout ),
    .A2(\__uuf__._0461_ ),
    .B1(\__uuf__.shifter.shiftreg[23] ),
    .B2(\__uuf__._0460_ ),
    .X(\__uuf__._0109_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1324_ 
  (
    .A1(\__BoundaryScanRegister_input_55__.dout ),
    .A2(\__uuf__._0461_ ),
    .B1(\__uuf__.shifter.shiftreg[24] ),
    .B2(\__uuf__._0460_ ),
    .X(\__uuf__._0110_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1325_ 
  (
    .A1(\__BoundaryScanRegister_input_56__.dout ),
    .A2(\__uuf__._0461_ ),
    .B1(\__uuf__.shifter.shiftreg[25] ),
    .B2(\__uuf__._0460_ ),
    .X(\__uuf__._0111_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1326_ 
  (
    .A(\__uuf__._0457_ ),
    .X(\__uuf__._0462_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1327_ 
  (
    .A1(\__BoundaryScanRegister_input_57__.dout ),
    .A2(\__uuf__._0461_ ),
    .B1(\__uuf__.shifter.shiftreg[26] ),
    .B2(\__uuf__._0462_ ),
    .X(\__uuf__._0112_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1328_ 
  (
    .A1(\__BoundaryScanRegister_input_58__.dout ),
    .A2(\__uuf__._0461_ ),
    .B1(\__uuf__.shifter.shiftreg[27] ),
    .B2(\__uuf__._0462_ ),
    .X(\__uuf__._0113_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1329_ 
  (
    .A(\__uuf__._0807_ ),
    .X(\__uuf__._0463_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1330_ 
  (
    .A1(\__BoundaryScanRegister_input_59__.dout ),
    .A2(\__uuf__._0463_ ),
    .B1(\__uuf__.shifter.shiftreg[28] ),
    .B2(\__uuf__._0462_ ),
    .X(\__uuf__._0114_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1331_ 
  (
    .A1(\__BoundaryScanRegister_input_60__.dout ),
    .A2(\__uuf__._0463_ ),
    .B1(\__uuf__.shifter.shiftreg[29] ),
    .B2(\__uuf__._0462_ ),
    .X(\__uuf__._0115_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1332_ 
  (
    .A1(\__BoundaryScanRegister_input_61__.dout ),
    .A2(\__uuf__._0463_ ),
    .B1(\__uuf__.shifter.shiftreg[30] ),
    .B2(\__uuf__._0462_ ),
    .X(\__uuf__._0116_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1333_ 
  (
    .A(\__uuf__._0457_ ),
    .X(\__uuf__._0464_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1334_ 
  (
    .A1(\__BoundaryScanRegister_input_62__.dout ),
    .A2(\__uuf__._0463_ ),
    .B1(\__uuf__.shifter.shiftreg[31] ),
    .B2(\__uuf__._0464_ ),
    .X(\__uuf__._0118_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1335_ 
  (
    .A(\__uuf__._0865_ ),
    .X(\__uuf__._0465_ )
  );


  sky130_fd_sc_hd__and2_4
  \__uuf__._1336_ 
  (
    .A(\__BoundaryScanRegister_input_63__.dout ),
    .B(\__uuf__._0788_ ),
    .X(\__uuf__._0466_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1337_ 
  (
    .A(\__uuf__._0466_ ),
    .X(\__uuf__._0467_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1338_ 
  (
    .A(\__uuf__._0467_ ),
    .X(\__uuf__._0154_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1339_ 
  (
    .A1(\__uuf__.shifter.shiftreg[32] ),
    .A2(\__uuf__._0465_ ),
    .B1(\__uuf__._0154_ ),
    .X(\__uuf__._0119_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1340_ 
  (
    .A1(\__uuf__.shifter.shiftreg[33] ),
    .A2(\__uuf__._0465_ ),
    .B1(\__uuf__._0154_ ),
    .X(\__uuf__._0120_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1341_ 
  (
    .A1(\__uuf__.shifter.shiftreg[34] ),
    .A2(\__uuf__._0465_ ),
    .B1(\__uuf__._0154_ ),
    .X(\__uuf__._0121_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1342_ 
  (
    .A1(\__uuf__.shifter.shiftreg[35] ),
    .A2(\__uuf__._0465_ ),
    .B1(\__uuf__._0154_ ),
    .X(\__uuf__._0122_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1343_ 
  (
    .A(\__uuf__._0467_ ),
    .X(\__uuf__._0468_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1344_ 
  (
    .A(\__uuf__._0468_ ),
    .X(\__uuf__._0469_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1345_ 
  (
    .A1(\__uuf__.shifter.shiftreg[36] ),
    .A2(\__uuf__._0465_ ),
    .B1(\__uuf__._0469_ ),
    .X(\__uuf__._0123_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1346_ 
  (
    .A(\__uuf__._0860_ ),
    .X(\__uuf__._0470_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1347_ 
  (
    .A(\__uuf__._0470_ ),
    .X(\__uuf__._0471_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1348_ 
  (
    .A1(\__uuf__.shifter.shiftreg[37] ),
    .A2(\__uuf__._0471_ ),
    .B1(\__uuf__._0469_ ),
    .X(\__uuf__._0124_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1349_ 
  (
    .A1(\__uuf__.shifter.shiftreg[38] ),
    .A2(\__uuf__._0471_ ),
    .B1(\__uuf__._0469_ ),
    .X(\__uuf__._0125_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1350_ 
  (
    .A1(\__uuf__.shifter.shiftreg[39] ),
    .A2(\__uuf__._0471_ ),
    .B1(\__uuf__._0469_ ),
    .X(\__uuf__._0126_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1351_ 
  (
    .A1(\__uuf__.shifter.shiftreg[40] ),
    .A2(\__uuf__._0471_ ),
    .B1(\__uuf__._0469_ ),
    .X(\__uuf__._0127_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1352_ 
  (
    .A(\__uuf__._0468_ ),
    .X(\__uuf__._0472_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1353_ 
  (
    .A1(\__uuf__.shifter.shiftreg[41] ),
    .A2(\__uuf__._0471_ ),
    .B1(\__uuf__._0472_ ),
    .X(\__uuf__._0129_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1354_ 
  (
    .A(\__uuf__._0470_ ),
    .X(\__uuf__._0473_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1355_ 
  (
    .A1(\__uuf__.shifter.shiftreg[42] ),
    .A2(\__uuf__._0473_ ),
    .B1(\__uuf__._0472_ ),
    .X(\__uuf__._0130_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1356_ 
  (
    .A1(\__uuf__.shifter.shiftreg[43] ),
    .A2(\__uuf__._0473_ ),
    .B1(\__uuf__._0472_ ),
    .X(\__uuf__._0131_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1357_ 
  (
    .A1(\__uuf__.shifter.shiftreg[44] ),
    .A2(\__uuf__._0473_ ),
    .B1(\__uuf__._0472_ ),
    .X(\__uuf__._0132_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1358_ 
  (
    .A1(\__uuf__.shifter.shiftreg[45] ),
    .A2(\__uuf__._0473_ ),
    .B1(\__uuf__._0472_ ),
    .X(\__uuf__._0133_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1359_ 
  (
    .A(\__uuf__._0467_ ),
    .X(\__uuf__._0474_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1360_ 
  (
    .A1(\__uuf__.shifter.shiftreg[46] ),
    .A2(\__uuf__._0473_ ),
    .B1(\__uuf__._0474_ ),
    .X(\__uuf__._0134_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1361_ 
  (
    .A(\__uuf__._0470_ ),
    .X(\__uuf__._0475_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1362_ 
  (
    .A1(\__uuf__.shifter.shiftreg[47] ),
    .A2(\__uuf__._0475_ ),
    .B1(\__uuf__._0474_ ),
    .X(\__uuf__._0135_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1363_ 
  (
    .A1(\__uuf__.shifter.shiftreg[48] ),
    .A2(\__uuf__._0475_ ),
    .B1(\__uuf__._0474_ ),
    .X(\__uuf__._0136_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1364_ 
  (
    .A1(\__uuf__.shifter.shiftreg[49] ),
    .A2(\__uuf__._0475_ ),
    .B1(\__uuf__._0474_ ),
    .X(\__uuf__._0137_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1365_ 
  (
    .A1(\__uuf__.shifter.shiftreg[50] ),
    .A2(\__uuf__._0475_ ),
    .B1(\__uuf__._0474_ ),
    .X(\__uuf__._0138_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1366_ 
  (
    .A(\__uuf__._0467_ ),
    .X(\__uuf__._0476_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1367_ 
  (
    .A1(\__uuf__.shifter.shiftreg[51] ),
    .A2(\__uuf__._0475_ ),
    .B1(\__uuf__._0476_ ),
    .X(\__uuf__._0140_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1368_ 
  (
    .A(\__uuf__._0470_ ),
    .X(\__uuf__._0477_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1369_ 
  (
    .A1(\__uuf__.shifter.shiftreg[52] ),
    .A2(\__uuf__._0477_ ),
    .B1(\__uuf__._0476_ ),
    .X(\__uuf__._0141_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1370_ 
  (
    .A1(\__uuf__.shifter.shiftreg[53] ),
    .A2(\__uuf__._0477_ ),
    .B1(\__uuf__._0476_ ),
    .X(\__uuf__._0142_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1371_ 
  (
    .A1(\__uuf__.shifter.shiftreg[54] ),
    .A2(\__uuf__._0477_ ),
    .B1(\__uuf__._0476_ ),
    .X(\__uuf__._0143_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1372_ 
  (
    .A1(\__uuf__.shifter.shiftreg[55] ),
    .A2(\__uuf__._0477_ ),
    .B1(\__uuf__._0476_ ),
    .X(\__uuf__._0144_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1373_ 
  (
    .A(\__uuf__._0467_ ),
    .X(\__uuf__._0478_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1374_ 
  (
    .A1(\__uuf__.shifter.shiftreg[56] ),
    .A2(\__uuf__._0477_ ),
    .B1(\__uuf__._0478_ ),
    .X(\__uuf__._0145_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1375_ 
  (
    .A(\__uuf__._0470_ ),
    .X(\__uuf__._0479_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1376_ 
  (
    .A1(\__uuf__.shifter.shiftreg[57] ),
    .A2(\__uuf__._0479_ ),
    .B1(\__uuf__._0478_ ),
    .X(\__uuf__._0146_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1377_ 
  (
    .A1(\__uuf__.shifter.shiftreg[58] ),
    .A2(\__uuf__._0479_ ),
    .B1(\__uuf__._0478_ ),
    .X(\__uuf__._0147_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1378_ 
  (
    .A1(\__uuf__.shifter.shiftreg[59] ),
    .A2(\__uuf__._0479_ ),
    .B1(\__uuf__._0478_ ),
    .X(\__uuf__._0148_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1379_ 
  (
    .A1(\__uuf__.shifter.shiftreg[60] ),
    .A2(\__uuf__._0479_ ),
    .B1(\__uuf__._0478_ ),
    .X(\__uuf__._0149_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1380_ 
  (
    .A1(\__uuf__.shifter.shiftreg[61] ),
    .A2(\__uuf__._0479_ ),
    .B1(\__uuf__._0468_ ),
    .X(\__uuf__._0151_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1381_ 
  (
    .A1(\__uuf__.shifter.shiftreg[62] ),
    .A2(\__uuf__._0447_ ),
    .B1(\__uuf__._0468_ ),
    .X(\__uuf__._0152_ )
  );


  sky130_fd_sc_hd__a21o_4
  \__uuf__._1382_ 
  (
    .A1(\__uuf__.shifter.shiftreg[63] ),
    .A2(\__uuf__._0447_ ),
    .B1(\__uuf__._0468_ ),
    .X(\__uuf__._0153_ )
  );


  sky130_fd_sc_hd__and2_4
  \__uuf__._1383_ 
  (
    .A(\__uuf__.shifter.shiftreg[0] ),
    .B(\__uuf__._0447_ ),
    .X(\__uuf__._0094_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1384_ 
  (
    .A(\__uuf__._0083_ ),
    .Y(\__uuf__._0480_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1385_ 
  (
    .A(\__uuf__.multiplier.pp[31] ),
    .Y(\__uuf__._0481_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1386_ 
  (
    .A(\__uuf__.multiplier.y ),
    .Y(\__uuf__._0482_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1387_ 
  (
    .A(\__uuf__._0482_ ),
    .X(\__uuf__._0483_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1388_ 
  (
    .A(\__BoundaryScanRegister_input_30__.dout ),
    .Y(\__uuf__._0484_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1389_ 
  (
    .A1(\__uuf__._0480_ ),
    .A2(\__uuf__._0481_ ),
    .B1(\__uuf__._0483_ ),
    .B2(\__uuf__._0484_ ),
    .X(\__uuf__._0485_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1390_ 
  (
    .A1(\__uuf__._0480_ ),
    .A2(\__uuf__._0481_ ),
    .B1(\__uuf__._0464_ ),
    .C1(\__uuf__._0485_ ),
    .X(\__uuf__._0486_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1391_ 
  (
    .A(\__uuf__._0486_ ),
    .Y(\__uuf__._0081_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1392_ 
  (
    .A(\__uuf__._0482_ ),
    .X(\__uuf__._0487_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1393_ 
  (
    .A(\__uuf__._0487_ ),
    .X(\__uuf__._0488_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1394_ 
  (
    .A1_N(\__uuf__._0480_ ),
    .A2_N(\__uuf__._0481_ ),
    .B1(\__uuf__._0480_ ),
    .B2(\__uuf__._0481_ ),
    .X(\__uuf__._0489_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1395_ 
  (
    .A(\__uuf__._0488_ ),
    .B(\__uuf__._0484_ ),
    .C(\__uuf__._0489_ ),
    .X(\__uuf__._0490_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1396_ 
  (
    .A(\__uuf__._0482_ ),
    .X(\__uuf__._0491_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1397_ 
  (
    .A(\__uuf__._0491_ ),
    .X(\__uuf__._0492_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1398_ 
  (
    .A1(\__uuf__._0492_ ),
    .A2(\__uuf__._0484_ ),
    .B1(\__uuf__._0489_ ),
    .Y(\__uuf__._0493_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1399_ 
  (
    .A(\__uuf__._0463_ ),
    .B(\__uuf__._0490_ ),
    .C(\__uuf__._0493_ ),
    .X(\__uuf__._0082_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1400_ 
  (
    .A(\__uuf__._0080_ ),
    .Y(\__uuf__._0494_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1401_ 
  (
    .A(\__uuf__.multiplier.pp[30] ),
    .Y(\__uuf__._0495_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1402_ 
  (
    .A(\__BoundaryScanRegister_input_29__.dout ),
    .Y(\__uuf__._0496_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1403_ 
  (
    .A1(\__uuf__._0494_ ),
    .A2(\__uuf__._0495_ ),
    .B1(\__uuf__._0483_ ),
    .B2(\__uuf__._0496_ ),
    .X(\__uuf__._0497_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1404_ 
  (
    .A1(\__uuf__._0494_ ),
    .A2(\__uuf__._0495_ ),
    .B1(\__uuf__._0464_ ),
    .C1(\__uuf__._0497_ ),
    .X(\__uuf__._0498_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1405_ 
  (
    .A(\__uuf__._0498_ ),
    .Y(\__uuf__._0078_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1406_ 
  (
    .A(\__uuf__._0860_ ),
    .X(\__uuf__._0499_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1407_ 
  (
    .A(\__uuf__._0499_ ),
    .X(\__uuf__._0500_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1408_ 
  (
    .A1_N(\__uuf__._0494_ ),
    .A2_N(\__uuf__._0495_ ),
    .B1(\__uuf__._0494_ ),
    .B2(\__uuf__._0495_ ),
    .X(\__uuf__._0501_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1409_ 
  (
    .A(\__uuf__._0488_ ),
    .B(\__uuf__._0496_ ),
    .C(\__uuf__._0501_ ),
    .X(\__uuf__._0502_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1410_ 
  (
    .A1(\__uuf__._0492_ ),
    .A2(\__uuf__._0496_ ),
    .B1(\__uuf__._0501_ ),
    .Y(\__uuf__._0503_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1411_ 
  (
    .A(\__uuf__._0500_ ),
    .B(\__uuf__._0502_ ),
    .C(\__uuf__._0503_ ),
    .X(\__uuf__._0079_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1412_ 
  (
    .A(\__uuf__._0077_ ),
    .Y(\__uuf__._0504_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1413_ 
  (
    .A(\__uuf__.multiplier.pp[29] ),
    .Y(\__uuf__._0505_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1414_ 
  (
    .A(\__BoundaryScanRegister_input_28__.dout ),
    .Y(\__uuf__._0506_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1415_ 
  (
    .A1(\__uuf__._0504_ ),
    .A2(\__uuf__._0505_ ),
    .B1(\__uuf__._0483_ ),
    .B2(\__uuf__._0506_ ),
    .X(\__uuf__._0507_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1416_ 
  (
    .A1(\__uuf__._0504_ ),
    .A2(\__uuf__._0505_ ),
    .B1(\__uuf__._0464_ ),
    .C1(\__uuf__._0507_ ),
    .X(\__uuf__._0508_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1417_ 
  (
    .A(\__uuf__._0508_ ),
    .Y(\__uuf__._0075_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1418_ 
  (
    .A1_N(\__uuf__._0504_ ),
    .A2_N(\__uuf__._0505_ ),
    .B1(\__uuf__._0504_ ),
    .B2(\__uuf__._0505_ ),
    .X(\__uuf__._0509_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1419_ 
  (
    .A(\__uuf__._0488_ ),
    .B(\__uuf__._0506_ ),
    .C(\__uuf__._0509_ ),
    .X(\__uuf__._0510_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1420_ 
  (
    .A1(\__uuf__._0492_ ),
    .A2(\__uuf__._0506_ ),
    .B1(\__uuf__._0509_ ),
    .Y(\__uuf__._0511_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1421_ 
  (
    .A(\__uuf__._0500_ ),
    .B(\__uuf__._0510_ ),
    .C(\__uuf__._0511_ ),
    .X(\__uuf__._0076_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1422_ 
  (
    .A(\__uuf__._0074_ ),
    .Y(\__uuf__._0512_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1423_ 
  (
    .A(\__uuf__.multiplier.pp[28] ),
    .Y(\__uuf__._0513_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1424_ 
  (
    .A(\__uuf__._0482_ ),
    .X(\__uuf__._0514_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1425_ 
  (
    .A(\__uuf__._0514_ ),
    .X(\__uuf__._0515_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1426_ 
  (
    .A(\__BoundaryScanRegister_input_27__.dout ),
    .Y(\__uuf__._0516_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1427_ 
  (
    .A1(\__uuf__._0512_ ),
    .A2(\__uuf__._0513_ ),
    .B1(\__uuf__._0515_ ),
    .B2(\__uuf__._0516_ ),
    .X(\__uuf__._0517_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1428_ 
  (
    .A1(\__uuf__._0512_ ),
    .A2(\__uuf__._0513_ ),
    .B1(\__uuf__._0464_ ),
    .C1(\__uuf__._0517_ ),
    .X(\__uuf__._0518_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1429_ 
  (
    .A(\__uuf__._0518_ ),
    .Y(\__uuf__._0072_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1430_ 
  (
    .A1_N(\__uuf__._0512_ ),
    .A2_N(\__uuf__._0513_ ),
    .B1(\__uuf__._0512_ ),
    .B2(\__uuf__._0513_ ),
    .X(\__uuf__._0519_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1431_ 
  (
    .A(\__uuf__._0488_ ),
    .B(\__uuf__._0516_ ),
    .C(\__uuf__._0519_ ),
    .X(\__uuf__._0520_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1432_ 
  (
    .A1(\__uuf__._0492_ ),
    .A2(\__uuf__._0516_ ),
    .B1(\__uuf__._0519_ ),
    .Y(\__uuf__._0521_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1433_ 
  (
    .A(\__uuf__._0500_ ),
    .B(\__uuf__._0520_ ),
    .C(\__uuf__._0521_ ),
    .X(\__uuf__._0073_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1434_ 
  (
    .A(\__uuf__._0071_ ),
    .Y(\__uuf__._0522_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1435_ 
  (
    .A(\__uuf__.multiplier.pp[27] ),
    .Y(\__uuf__._0523_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1436_ 
  (
    .A(\__uuf__._0457_ ),
    .X(\__uuf__._0524_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1437_ 
  (
    .A(\__BoundaryScanRegister_input_26__.dout ),
    .Y(\__uuf__._0525_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1438_ 
  (
    .A1(\__uuf__._0522_ ),
    .A2(\__uuf__._0523_ ),
    .B1(\__uuf__._0515_ ),
    .B2(\__uuf__._0525_ ),
    .X(\__uuf__._0526_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1439_ 
  (
    .A1(\__uuf__._0522_ ),
    .A2(\__uuf__._0523_ ),
    .B1(\__uuf__._0524_ ),
    .C1(\__uuf__._0526_ ),
    .X(\__uuf__._0527_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1440_ 
  (
    .A(\__uuf__._0527_ ),
    .Y(\__uuf__._0069_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1441_ 
  (
    .A(\__uuf__._0482_ ),
    .X(\__uuf__._0528_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1442_ 
  (
    .A(\__uuf__._0528_ ),
    .X(\__uuf__._0529_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1443_ 
  (
    .A1_N(\__uuf__._0522_ ),
    .A2_N(\__uuf__._0523_ ),
    .B1(\__uuf__._0522_ ),
    .B2(\__uuf__._0523_ ),
    .X(\__uuf__._0530_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1444_ 
  (
    .A(\__uuf__._0529_ ),
    .B(\__uuf__._0525_ ),
    .C(\__uuf__._0530_ ),
    .X(\__uuf__._0531_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1445_ 
  (
    .A1(\__uuf__._0492_ ),
    .A2(\__uuf__._0525_ ),
    .B1(\__uuf__._0530_ ),
    .Y(\__uuf__._0532_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1446_ 
  (
    .A(\__uuf__._0500_ ),
    .B(\__uuf__._0531_ ),
    .C(\__uuf__._0532_ ),
    .X(\__uuf__._0070_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1447_ 
  (
    .A(\__uuf__._0068_ ),
    .Y(\__uuf__._0533_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1448_ 
  (
    .A(\__uuf__.multiplier.pp[26] ),
    .Y(\__uuf__._0534_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1449_ 
  (
    .A(\__BoundaryScanRegister_input_25__.dout ),
    .Y(\__uuf__._0535_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1450_ 
  (
    .A1(\__uuf__._0533_ ),
    .A2(\__uuf__._0534_ ),
    .B1(\__uuf__._0515_ ),
    .B2(\__uuf__._0535_ ),
    .X(\__uuf__._0536_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1451_ 
  (
    .A1(\__uuf__._0533_ ),
    .A2(\__uuf__._0534_ ),
    .B1(\__uuf__._0524_ ),
    .C1(\__uuf__._0536_ ),
    .X(\__uuf__._0537_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1452_ 
  (
    .A(\__uuf__._0537_ ),
    .Y(\__uuf__._0066_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1453_ 
  (
    .A1_N(\__uuf__._0533_ ),
    .A2_N(\__uuf__._0534_ ),
    .B1(\__uuf__._0533_ ),
    .B2(\__uuf__._0534_ ),
    .X(\__uuf__._0538_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1454_ 
  (
    .A(\__uuf__._0529_ ),
    .B(\__uuf__._0535_ ),
    .C(\__uuf__._0538_ ),
    .X(\__uuf__._0539_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1455_ 
  (
    .A(\__uuf__._0491_ ),
    .X(\__uuf__._0540_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1456_ 
  (
    .A1(\__uuf__._0540_ ),
    .A2(\__uuf__._0535_ ),
    .B1(\__uuf__._0538_ ),
    .Y(\__uuf__._0541_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1457_ 
  (
    .A(\__uuf__._0500_ ),
    .B(\__uuf__._0539_ ),
    .C(\__uuf__._0541_ ),
    .X(\__uuf__._0067_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1458_ 
  (
    .A(\__uuf__._0065_ ),
    .Y(\__uuf__._0542_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1459_ 
  (
    .A(\__uuf__.multiplier.pp[25] ),
    .Y(\__uuf__._0543_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1460_ 
  (
    .A(\__BoundaryScanRegister_input_24__.dout ),
    .Y(\__uuf__._0544_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1461_ 
  (
    .A1(\__uuf__._0542_ ),
    .A2(\__uuf__._0543_ ),
    .B1(\__uuf__._0515_ ),
    .B2(\__uuf__._0544_ ),
    .X(\__uuf__._0545_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1462_ 
  (
    .A1(\__uuf__._0542_ ),
    .A2(\__uuf__._0543_ ),
    .B1(\__uuf__._0524_ ),
    .C1(\__uuf__._0545_ ),
    .X(\__uuf__._0546_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1463_ 
  (
    .A(\__uuf__._0546_ ),
    .Y(\__uuf__._0063_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1464_ 
  (
    .A(\__uuf__._0499_ ),
    .X(\__uuf__._0547_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1465_ 
  (
    .A1_N(\__uuf__._0542_ ),
    .A2_N(\__uuf__._0543_ ),
    .B1(\__uuf__._0542_ ),
    .B2(\__uuf__._0543_ ),
    .X(\__uuf__._0548_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1466_ 
  (
    .A(\__uuf__._0529_ ),
    .B(\__uuf__._0544_ ),
    .C(\__uuf__._0548_ ),
    .X(\__uuf__._0549_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1467_ 
  (
    .A1(\__uuf__._0540_ ),
    .A2(\__uuf__._0544_ ),
    .B1(\__uuf__._0548_ ),
    .Y(\__uuf__._0550_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1468_ 
  (
    .A(\__uuf__._0547_ ),
    .B(\__uuf__._0549_ ),
    .C(\__uuf__._0550_ ),
    .X(\__uuf__._0064_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1469_ 
  (
    .A(\__uuf__._0062_ ),
    .Y(\__uuf__._0551_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1470_ 
  (
    .A(\__uuf__.multiplier.pp[24] ),
    .Y(\__uuf__._0552_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1471_ 
  (
    .A(\__BoundaryScanRegister_input_23__.dout ),
    .Y(\__uuf__._0553_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1472_ 
  (
    .A1(\__uuf__._0551_ ),
    .A2(\__uuf__._0552_ ),
    .B1(\__uuf__._0515_ ),
    .B2(\__uuf__._0553_ ),
    .X(\__uuf__._0554_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1473_ 
  (
    .A1(\__uuf__._0551_ ),
    .A2(\__uuf__._0552_ ),
    .B1(\__uuf__._0524_ ),
    .C1(\__uuf__._0554_ ),
    .X(\__uuf__._0555_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1474_ 
  (
    .A(\__uuf__._0555_ ),
    .Y(\__uuf__._0060_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1475_ 
  (
    .A1_N(\__uuf__._0551_ ),
    .A2_N(\__uuf__._0552_ ),
    .B1(\__uuf__._0551_ ),
    .B2(\__uuf__._0552_ ),
    .X(\__uuf__._0556_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1476_ 
  (
    .A(\__uuf__._0529_ ),
    .B(\__uuf__._0553_ ),
    .C(\__uuf__._0556_ ),
    .X(\__uuf__._0557_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1477_ 
  (
    .A1(\__uuf__._0540_ ),
    .A2(\__uuf__._0553_ ),
    .B1(\__uuf__._0556_ ),
    .Y(\__uuf__._0558_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1478_ 
  (
    .A(\__uuf__._0547_ ),
    .B(\__uuf__._0557_ ),
    .C(\__uuf__._0558_ ),
    .X(\__uuf__._0061_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1479_ 
  (
    .A(\__uuf__._0059_ ),
    .Y(\__uuf__._0559_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1480_ 
  (
    .A(\__uuf__.multiplier.pp[23] ),
    .Y(\__uuf__._0560_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1481_ 
  (
    .A(\__uuf__._0514_ ),
    .X(\__uuf__._0561_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1482_ 
  (
    .A(\__BoundaryScanRegister_input_22__.dout ),
    .Y(\__uuf__._0562_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1483_ 
  (
    .A1(\__uuf__._0559_ ),
    .A2(\__uuf__._0560_ ),
    .B1(\__uuf__._0561_ ),
    .B2(\__uuf__._0562_ ),
    .X(\__uuf__._0563_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1484_ 
  (
    .A1(\__uuf__._0559_ ),
    .A2(\__uuf__._0560_ ),
    .B1(\__uuf__._0524_ ),
    .C1(\__uuf__._0563_ ),
    .X(\__uuf__._0564_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1485_ 
  (
    .A(\__uuf__._0564_ ),
    .Y(\__uuf__._0057_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1486_ 
  (
    .A1_N(\__uuf__._0559_ ),
    .A2_N(\__uuf__._0560_ ),
    .B1(\__uuf__._0559_ ),
    .B2(\__uuf__._0560_ ),
    .X(\__uuf__._0565_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1487_ 
  (
    .A(\__uuf__._0529_ ),
    .B(\__uuf__._0562_ ),
    .C(\__uuf__._0565_ ),
    .X(\__uuf__._0566_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1488_ 
  (
    .A1(\__uuf__._0540_ ),
    .A2(\__uuf__._0562_ ),
    .B1(\__uuf__._0565_ ),
    .Y(\__uuf__._0567_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1489_ 
  (
    .A(\__uuf__._0547_ ),
    .B(\__uuf__._0566_ ),
    .C(\__uuf__._0567_ ),
    .X(\__uuf__._0058_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1490_ 
  (
    .A(\__uuf__._0056_ ),
    .Y(\__uuf__._0568_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1491_ 
  (
    .A(\__uuf__.multiplier.pp[22] ),
    .Y(\__uuf__._0569_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1492_ 
  (
    .A(\__uuf__._0448_ ),
    .X(\__uuf__._0570_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1493_ 
  (
    .A(\__BoundaryScanRegister_input_21__.dout ),
    .Y(\__uuf__._0571_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1494_ 
  (
    .A1(\__uuf__._0568_ ),
    .A2(\__uuf__._0569_ ),
    .B1(\__uuf__._0561_ ),
    .B2(\__uuf__._0571_ ),
    .X(\__uuf__._0572_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1495_ 
  (
    .A1(\__uuf__._0568_ ),
    .A2(\__uuf__._0569_ ),
    .B1(\__uuf__._0570_ ),
    .C1(\__uuf__._0572_ ),
    .X(\__uuf__._0573_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1496_ 
  (
    .A(\__uuf__._0573_ ),
    .Y(\__uuf__._0054_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1497_ 
  (
    .A(\__uuf__._0487_ ),
    .X(\__uuf__._0574_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1498_ 
  (
    .A1_N(\__uuf__._0568_ ),
    .A2_N(\__uuf__._0569_ ),
    .B1(\__uuf__._0568_ ),
    .B2(\__uuf__._0569_ ),
    .X(\__uuf__._0575_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1499_ 
  (
    .A(\__uuf__._0574_ ),
    .B(\__uuf__._0571_ ),
    .C(\__uuf__._0575_ ),
    .X(\__uuf__._0576_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1500_ 
  (
    .A1(\__uuf__._0540_ ),
    .A2(\__uuf__._0571_ ),
    .B1(\__uuf__._0575_ ),
    .Y(\__uuf__._0577_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1501_ 
  (
    .A(\__uuf__._0547_ ),
    .B(\__uuf__._0576_ ),
    .C(\__uuf__._0577_ ),
    .X(\__uuf__._0055_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1502_ 
  (
    .A(\__uuf__._0053_ ),
    .Y(\__uuf__._0578_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1503_ 
  (
    .A(\__uuf__.multiplier.pp[21] ),
    .Y(\__uuf__._0579_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1504_ 
  (
    .A(\__BoundaryScanRegister_input_20__.dout ),
    .Y(\__uuf__._0580_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1505_ 
  (
    .A1(\__uuf__._0578_ ),
    .A2(\__uuf__._0579_ ),
    .B1(\__uuf__._0561_ ),
    .B2(\__uuf__._0580_ ),
    .X(\__uuf__._0581_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1506_ 
  (
    .A1(\__uuf__._0578_ ),
    .A2(\__uuf__._0579_ ),
    .B1(\__uuf__._0570_ ),
    .C1(\__uuf__._0581_ ),
    .X(\__uuf__._0582_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1507_ 
  (
    .A(\__uuf__._0582_ ),
    .Y(\__uuf__._0051_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1508_ 
  (
    .A1_N(\__uuf__._0578_ ),
    .A2_N(\__uuf__._0579_ ),
    .B1(\__uuf__._0578_ ),
    .B2(\__uuf__._0579_ ),
    .X(\__uuf__._0583_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1509_ 
  (
    .A(\__uuf__._0574_ ),
    .B(\__uuf__._0580_ ),
    .C(\__uuf__._0583_ ),
    .X(\__uuf__._0584_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1510_ 
  (
    .A(\__uuf__._0528_ ),
    .X(\__uuf__._0585_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1511_ 
  (
    .A1(\__uuf__._0585_ ),
    .A2(\__uuf__._0580_ ),
    .B1(\__uuf__._0583_ ),
    .Y(\__uuf__._0586_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1512_ 
  (
    .A(\__uuf__._0547_ ),
    .B(\__uuf__._0584_ ),
    .C(\__uuf__._0586_ ),
    .X(\__uuf__._0052_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1513_ 
  (
    .A(\__uuf__._0050_ ),
    .Y(\__uuf__._0587_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1514_ 
  (
    .A(\__uuf__.multiplier.pp[20] ),
    .Y(\__uuf__._0588_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1515_ 
  (
    .A(\__BoundaryScanRegister_input_19__.dout ),
    .Y(\__uuf__._0589_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1516_ 
  (
    .A1(\__uuf__._0587_ ),
    .A2(\__uuf__._0588_ ),
    .B1(\__uuf__._0561_ ),
    .B2(\__uuf__._0589_ ),
    .X(\__uuf__._0590_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1517_ 
  (
    .A1(\__uuf__._0587_ ),
    .A2(\__uuf__._0588_ ),
    .B1(\__uuf__._0570_ ),
    .C1(\__uuf__._0590_ ),
    .X(\__uuf__._0591_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1518_ 
  (
    .A(\__uuf__._0591_ ),
    .Y(\__uuf__._0048_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1519_ 
  (
    .A(\__uuf__._0499_ ),
    .X(\__uuf__._0592_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1520_ 
  (
    .A1_N(\__uuf__._0587_ ),
    .A2_N(\__uuf__._0588_ ),
    .B1(\__uuf__._0587_ ),
    .B2(\__uuf__._0588_ ),
    .X(\__uuf__._0593_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1521_ 
  (
    .A(\__uuf__._0574_ ),
    .B(\__uuf__._0589_ ),
    .C(\__uuf__._0593_ ),
    .X(\__uuf__._0594_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1522_ 
  (
    .A1(\__uuf__._0585_ ),
    .A2(\__uuf__._0589_ ),
    .B1(\__uuf__._0593_ ),
    .Y(\__uuf__._0595_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1523_ 
  (
    .A(\__uuf__._0592_ ),
    .B(\__uuf__._0594_ ),
    .C(\__uuf__._0595_ ),
    .X(\__uuf__._0049_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1524_ 
  (
    .A(\__uuf__._0047_ ),
    .Y(\__uuf__._0596_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1525_ 
  (
    .A(\__uuf__.multiplier.pp[19] ),
    .Y(\__uuf__._0597_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1526_ 
  (
    .A(\__BoundaryScanRegister_input_18__.dout ),
    .Y(\__uuf__._0598_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1527_ 
  (
    .A1(\__uuf__._0596_ ),
    .A2(\__uuf__._0597_ ),
    .B1(\__uuf__._0561_ ),
    .B2(\__uuf__._0598_ ),
    .X(\__uuf__._0599_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1528_ 
  (
    .A1(\__uuf__._0596_ ),
    .A2(\__uuf__._0597_ ),
    .B1(\__uuf__._0570_ ),
    .C1(\__uuf__._0599_ ),
    .X(\__uuf__._0600_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1529_ 
  (
    .A(\__uuf__._0600_ ),
    .Y(\__uuf__._0045_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1530_ 
  (
    .A1_N(\__uuf__._0596_ ),
    .A2_N(\__uuf__._0597_ ),
    .B1(\__uuf__._0596_ ),
    .B2(\__uuf__._0597_ ),
    .X(\__uuf__._0601_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1531_ 
  (
    .A(\__uuf__._0574_ ),
    .B(\__uuf__._0598_ ),
    .C(\__uuf__._0601_ ),
    .X(\__uuf__._0602_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1532_ 
  (
    .A1(\__uuf__._0585_ ),
    .A2(\__uuf__._0598_ ),
    .B1(\__uuf__._0601_ ),
    .Y(\__uuf__._0603_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1533_ 
  (
    .A(\__uuf__._0592_ ),
    .B(\__uuf__._0602_ ),
    .C(\__uuf__._0603_ ),
    .X(\__uuf__._0046_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1534_ 
  (
    .A(\__uuf__._0044_ ),
    .Y(\__uuf__._0604_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1535_ 
  (
    .A(\__uuf__.multiplier.pp[18] ),
    .Y(\__uuf__._0605_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1536_ 
  (
    .A(\__uuf__._0514_ ),
    .X(\__uuf__._0606_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1537_ 
  (
    .A(\__BoundaryScanRegister_input_17__.dout ),
    .Y(\__uuf__._0607_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1538_ 
  (
    .A1(\__uuf__._0604_ ),
    .A2(\__uuf__._0605_ ),
    .B1(\__uuf__._0606_ ),
    .B2(\__uuf__._0607_ ),
    .X(\__uuf__._0608_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1539_ 
  (
    .A1(\__uuf__._0604_ ),
    .A2(\__uuf__._0605_ ),
    .B1(\__uuf__._0570_ ),
    .C1(\__uuf__._0608_ ),
    .X(\__uuf__._0609_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1540_ 
  (
    .A(\__uuf__._0609_ ),
    .Y(\__uuf__._0042_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1541_ 
  (
    .A1_N(\__uuf__._0604_ ),
    .A2_N(\__uuf__._0605_ ),
    .B1(\__uuf__._0604_ ),
    .B2(\__uuf__._0605_ ),
    .X(\__uuf__._0610_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1542_ 
  (
    .A(\__uuf__._0574_ ),
    .B(\__uuf__._0607_ ),
    .C(\__uuf__._0610_ ),
    .X(\__uuf__._0611_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1543_ 
  (
    .A1(\__uuf__._0585_ ),
    .A2(\__uuf__._0607_ ),
    .B1(\__uuf__._0610_ ),
    .Y(\__uuf__._0612_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1544_ 
  (
    .A(\__uuf__._0592_ ),
    .B(\__uuf__._0611_ ),
    .C(\__uuf__._0612_ ),
    .X(\__uuf__._0043_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1545_ 
  (
    .A(\__uuf__._0041_ ),
    .Y(\__uuf__._0613_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1546_ 
  (
    .A(\__uuf__.multiplier.pp[17] ),
    .Y(\__uuf__._0614_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1547_ 
  (
    .A(\__uuf__._0448_ ),
    .X(\__uuf__._0615_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1548_ 
  (
    .A(\__BoundaryScanRegister_input_16__.dout ),
    .Y(\__uuf__._0616_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1549_ 
  (
    .A1(\__uuf__._0613_ ),
    .A2(\__uuf__._0614_ ),
    .B1(\__uuf__._0606_ ),
    .B2(\__uuf__._0616_ ),
    .X(\__uuf__._0617_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1550_ 
  (
    .A1(\__uuf__._0613_ ),
    .A2(\__uuf__._0614_ ),
    .B1(\__uuf__._0615_ ),
    .C1(\__uuf__._0617_ ),
    .X(\__uuf__._0618_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1551_ 
  (
    .A(\__uuf__._0618_ ),
    .Y(\__uuf__._0039_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1552_ 
  (
    .A(\__uuf__._0487_ ),
    .X(\__uuf__._0619_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1553_ 
  (
    .A1_N(\__uuf__._0613_ ),
    .A2_N(\__uuf__._0614_ ),
    .B1(\__uuf__._0613_ ),
    .B2(\__uuf__._0614_ ),
    .X(\__uuf__._0620_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1554_ 
  (
    .A(\__uuf__._0619_ ),
    .B(\__uuf__._0616_ ),
    .C(\__uuf__._0620_ ),
    .X(\__uuf__._0621_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1555_ 
  (
    .A1(\__uuf__._0585_ ),
    .A2(\__uuf__._0616_ ),
    .B1(\__uuf__._0620_ ),
    .Y(\__uuf__._0622_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1556_ 
  (
    .A(\__uuf__._0592_ ),
    .B(\__uuf__._0621_ ),
    .C(\__uuf__._0622_ ),
    .X(\__uuf__._0040_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1557_ 
  (
    .A(\__uuf__._0038_ ),
    .Y(\__uuf__._0623_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1558_ 
  (
    .A(\__uuf__.multiplier.pp[16] ),
    .Y(\__uuf__._0624_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1559_ 
  (
    .A(\__BoundaryScanRegister_input_15__.dout ),
    .Y(\__uuf__._0625_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1560_ 
  (
    .A1(\__uuf__._0623_ ),
    .A2(\__uuf__._0624_ ),
    .B1(\__uuf__._0606_ ),
    .B2(\__uuf__._0625_ ),
    .X(\__uuf__._0626_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1561_ 
  (
    .A1(\__uuf__._0623_ ),
    .A2(\__uuf__._0624_ ),
    .B1(\__uuf__._0615_ ),
    .C1(\__uuf__._0626_ ),
    .X(\__uuf__._0627_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1562_ 
  (
    .A(\__uuf__._0627_ ),
    .Y(\__uuf__._0036_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1563_ 
  (
    .A1_N(\__uuf__._0623_ ),
    .A2_N(\__uuf__._0624_ ),
    .B1(\__uuf__._0623_ ),
    .B2(\__uuf__._0624_ ),
    .X(\__uuf__._0628_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1564_ 
  (
    .A(\__uuf__._0619_ ),
    .B(\__uuf__._0625_ ),
    .C(\__uuf__._0628_ ),
    .X(\__uuf__._0629_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1565_ 
  (
    .A(\__uuf__._0528_ ),
    .X(\__uuf__._0630_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1566_ 
  (
    .A1(\__uuf__._0630_ ),
    .A2(\__uuf__._0625_ ),
    .B1(\__uuf__._0628_ ),
    .Y(\__uuf__._0631_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1567_ 
  (
    .A(\__uuf__._0592_ ),
    .B(\__uuf__._0629_ ),
    .C(\__uuf__._0631_ ),
    .X(\__uuf__._0037_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1568_ 
  (
    .A(\__uuf__._0035_ ),
    .Y(\__uuf__._0632_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1569_ 
  (
    .A(\__uuf__.multiplier.pp[15] ),
    .Y(\__uuf__._0633_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1570_ 
  (
    .A(\__BoundaryScanRegister_input_14__.dout ),
    .Y(\__uuf__._0634_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1571_ 
  (
    .A1(\__uuf__._0632_ ),
    .A2(\__uuf__._0633_ ),
    .B1(\__uuf__._0606_ ),
    .B2(\__uuf__._0634_ ),
    .X(\__uuf__._0635_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1572_ 
  (
    .A1(\__uuf__._0632_ ),
    .A2(\__uuf__._0633_ ),
    .B1(\__uuf__._0615_ ),
    .C1(\__uuf__._0635_ ),
    .X(\__uuf__._0636_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1573_ 
  (
    .A(\__uuf__._0636_ ),
    .Y(\__uuf__._0033_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1574_ 
  (
    .A(\__uuf__._0499_ ),
    .X(\__uuf__._0637_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1575_ 
  (
    .A1_N(\__uuf__._0632_ ),
    .A2_N(\__uuf__._0633_ ),
    .B1(\__uuf__._0632_ ),
    .B2(\__uuf__._0633_ ),
    .X(\__uuf__._0638_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1576_ 
  (
    .A(\__uuf__._0619_ ),
    .B(\__uuf__._0634_ ),
    .C(\__uuf__._0638_ ),
    .X(\__uuf__._0639_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1577_ 
  (
    .A1(\__uuf__._0630_ ),
    .A2(\__uuf__._0634_ ),
    .B1(\__uuf__._0638_ ),
    .Y(\__uuf__._0640_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1578_ 
  (
    .A(\__uuf__._0637_ ),
    .B(\__uuf__._0639_ ),
    .C(\__uuf__._0640_ ),
    .X(\__uuf__._0034_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1579_ 
  (
    .A(\__uuf__._0032_ ),
    .Y(\__uuf__._0641_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1580_ 
  (
    .A(\__uuf__.multiplier.pp[14] ),
    .Y(\__uuf__._0642_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1581_ 
  (
    .A(\__BoundaryScanRegister_input_13__.dout ),
    .Y(\__uuf__._0643_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1582_ 
  (
    .A1(\__uuf__._0641_ ),
    .A2(\__uuf__._0642_ ),
    .B1(\__uuf__._0606_ ),
    .B2(\__uuf__._0643_ ),
    .X(\__uuf__._0644_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1583_ 
  (
    .A1(\__uuf__._0641_ ),
    .A2(\__uuf__._0642_ ),
    .B1(\__uuf__._0615_ ),
    .C1(\__uuf__._0644_ ),
    .X(\__uuf__._0645_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1584_ 
  (
    .A(\__uuf__._0645_ ),
    .Y(\__uuf__._0030_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1585_ 
  (
    .A1_N(\__uuf__._0641_ ),
    .A2_N(\__uuf__._0642_ ),
    .B1(\__uuf__._0641_ ),
    .B2(\__uuf__._0642_ ),
    .X(\__uuf__._0646_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1586_ 
  (
    .A(\__uuf__._0619_ ),
    .B(\__uuf__._0643_ ),
    .C(\__uuf__._0646_ ),
    .X(\__uuf__._0647_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1587_ 
  (
    .A1(\__uuf__._0630_ ),
    .A2(\__uuf__._0643_ ),
    .B1(\__uuf__._0646_ ),
    .Y(\__uuf__._0648_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1588_ 
  (
    .A(\__uuf__._0637_ ),
    .B(\__uuf__._0647_ ),
    .C(\__uuf__._0648_ ),
    .X(\__uuf__._0031_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1589_ 
  (
    .A(\__uuf__._0029_ ),
    .Y(\__uuf__._0649_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1590_ 
  (
    .A(\__uuf__.multiplier.pp[13] ),
    .Y(\__uuf__._0650_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1591_ 
  (
    .A(\__uuf__._0514_ ),
    .X(\__uuf__._0651_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1592_ 
  (
    .A(\__BoundaryScanRegister_input_12__.dout ),
    .Y(\__uuf__._0652_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1593_ 
  (
    .A1(\__uuf__._0649_ ),
    .A2(\__uuf__._0650_ ),
    .B1(\__uuf__._0651_ ),
    .B2(\__uuf__._0652_ ),
    .X(\__uuf__._0653_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1594_ 
  (
    .A1(\__uuf__._0649_ ),
    .A2(\__uuf__._0650_ ),
    .B1(\__uuf__._0615_ ),
    .C1(\__uuf__._0653_ ),
    .X(\__uuf__._0654_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1595_ 
  (
    .A(\__uuf__._0654_ ),
    .Y(\__uuf__._0027_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1596_ 
  (
    .A1_N(\__uuf__._0649_ ),
    .A2_N(\__uuf__._0650_ ),
    .B1(\__uuf__._0649_ ),
    .B2(\__uuf__._0650_ ),
    .X(\__uuf__._0655_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1597_ 
  (
    .A(\__uuf__._0619_ ),
    .B(\__uuf__._0652_ ),
    .C(\__uuf__._0655_ ),
    .X(\__uuf__._0656_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1598_ 
  (
    .A1(\__uuf__._0630_ ),
    .A2(\__uuf__._0652_ ),
    .B1(\__uuf__._0655_ ),
    .Y(\__uuf__._0657_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1599_ 
  (
    .A(\__uuf__._0637_ ),
    .B(\__uuf__._0656_ ),
    .C(\__uuf__._0657_ ),
    .X(\__uuf__._0028_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1600_ 
  (
    .A(\__uuf__._0026_ ),
    .Y(\__uuf__._0658_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1601_ 
  (
    .A(\__uuf__.multiplier.pp[12] ),
    .Y(\__uuf__._0659_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1602_ 
  (
    .A(\__uuf__._0448_ ),
    .X(\__uuf__._0660_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1603_ 
  (
    .A(\__BoundaryScanRegister_input_11__.dout ),
    .Y(\__uuf__._0661_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1604_ 
  (
    .A1(\__uuf__._0658_ ),
    .A2(\__uuf__._0659_ ),
    .B1(\__uuf__._0651_ ),
    .B2(\__uuf__._0661_ ),
    .X(\__uuf__._0662_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1605_ 
  (
    .A1(\__uuf__._0658_ ),
    .A2(\__uuf__._0659_ ),
    .B1(\__uuf__._0660_ ),
    .C1(\__uuf__._0662_ ),
    .X(\__uuf__._0663_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1606_ 
  (
    .A(\__uuf__._0663_ ),
    .Y(\__uuf__._0024_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1607_ 
  (
    .A(\__uuf__._0487_ ),
    .X(\__uuf__._0664_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1608_ 
  (
    .A1_N(\__uuf__._0658_ ),
    .A2_N(\__uuf__._0659_ ),
    .B1(\__uuf__._0658_ ),
    .B2(\__uuf__._0659_ ),
    .X(\__uuf__._0665_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1609_ 
  (
    .A(\__uuf__._0664_ ),
    .B(\__uuf__._0661_ ),
    .C(\__uuf__._0665_ ),
    .X(\__uuf__._0666_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1610_ 
  (
    .A1(\__uuf__._0630_ ),
    .A2(\__uuf__._0661_ ),
    .B1(\__uuf__._0665_ ),
    .Y(\__uuf__._0667_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1611_ 
  (
    .A(\__uuf__._0637_ ),
    .B(\__uuf__._0666_ ),
    .C(\__uuf__._0667_ ),
    .X(\__uuf__._0025_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1612_ 
  (
    .A(\__uuf__._0023_ ),
    .Y(\__uuf__._0668_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1613_ 
  (
    .A(\__uuf__.multiplier.pp[11] ),
    .Y(\__uuf__._0669_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1614_ 
  (
    .A(\__BoundaryScanRegister_input_10__.dout ),
    .Y(\__uuf__._0670_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1615_ 
  (
    .A1(\__uuf__._0668_ ),
    .A2(\__uuf__._0669_ ),
    .B1(\__uuf__._0651_ ),
    .B2(\__uuf__._0670_ ),
    .X(\__uuf__._0671_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1616_ 
  (
    .A1(\__uuf__._0668_ ),
    .A2(\__uuf__._0669_ ),
    .B1(\__uuf__._0660_ ),
    .C1(\__uuf__._0671_ ),
    .X(\__uuf__._0672_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1617_ 
  (
    .A(\__uuf__._0672_ ),
    .Y(\__uuf__._0021_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1618_ 
  (
    .A1_N(\__uuf__._0668_ ),
    .A2_N(\__uuf__._0669_ ),
    .B1(\__uuf__._0668_ ),
    .B2(\__uuf__._0669_ ),
    .X(\__uuf__._0673_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1619_ 
  (
    .A(\__uuf__._0664_ ),
    .B(\__uuf__._0670_ ),
    .C(\__uuf__._0673_ ),
    .X(\__uuf__._0674_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1620_ 
  (
    .A(\__uuf__._0528_ ),
    .X(\__uuf__._0675_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1621_ 
  (
    .A1(\__uuf__._0675_ ),
    .A2(\__uuf__._0670_ ),
    .B1(\__uuf__._0673_ ),
    .Y(\__uuf__._0676_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1622_ 
  (
    .A(\__uuf__._0637_ ),
    .B(\__uuf__._0674_ ),
    .C(\__uuf__._0676_ ),
    .X(\__uuf__._0022_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1623_ 
  (
    .A(\__uuf__._0020_ ),
    .Y(\__uuf__._0677_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1624_ 
  (
    .A(\__uuf__.multiplier.pp[10] ),
    .Y(\__uuf__._0678_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1625_ 
  (
    .A(\__BoundaryScanRegister_input_9__.dout ),
    .Y(\__uuf__._0679_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1626_ 
  (
    .A1(\__uuf__._0677_ ),
    .A2(\__uuf__._0678_ ),
    .B1(\__uuf__._0651_ ),
    .B2(\__uuf__._0679_ ),
    .X(\__uuf__._0680_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1627_ 
  (
    .A1(\__uuf__._0677_ ),
    .A2(\__uuf__._0678_ ),
    .B1(\__uuf__._0660_ ),
    .C1(\__uuf__._0680_ ),
    .X(\__uuf__._0681_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1628_ 
  (
    .A(\__uuf__._0681_ ),
    .Y(\__uuf__._0018_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1629_ 
  (
    .A(\__uuf__._0807_ ),
    .X(\__uuf__._0682_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1630_ 
  (
    .A1_N(\__uuf__._0677_ ),
    .A2_N(\__uuf__._0678_ ),
    .B1(\__uuf__._0677_ ),
    .B2(\__uuf__._0678_ ),
    .X(\__uuf__._0683_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1631_ 
  (
    .A(\__uuf__._0664_ ),
    .B(\__uuf__._0679_ ),
    .C(\__uuf__._0683_ ),
    .X(\__uuf__._0684_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1632_ 
  (
    .A1(\__uuf__._0675_ ),
    .A2(\__uuf__._0679_ ),
    .B1(\__uuf__._0683_ ),
    .Y(\__uuf__._0685_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1633_ 
  (
    .A(\__uuf__._0682_ ),
    .B(\__uuf__._0684_ ),
    .C(\__uuf__._0685_ ),
    .X(\__uuf__._0019_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1634_ 
  (
    .A(\__uuf__._0017_ ),
    .Y(\__uuf__._0686_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1635_ 
  (
    .A(\__uuf__.multiplier.pp[9] ),
    .Y(\__uuf__._0687_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1636_ 
  (
    .A(\__BoundaryScanRegister_input_8__.dout ),
    .Y(\__uuf__._0688_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1637_ 
  (
    .A1(\__uuf__._0686_ ),
    .A2(\__uuf__._0687_ ),
    .B1(\__uuf__._0651_ ),
    .B2(\__uuf__._0688_ ),
    .X(\__uuf__._0689_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1638_ 
  (
    .A1(\__uuf__._0686_ ),
    .A2(\__uuf__._0687_ ),
    .B1(\__uuf__._0660_ ),
    .C1(\__uuf__._0689_ ),
    .X(\__uuf__._0690_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1639_ 
  (
    .A(\__uuf__._0690_ ),
    .Y(\__uuf__._0015_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1640_ 
  (
    .A1_N(\__uuf__._0686_ ),
    .A2_N(\__uuf__._0687_ ),
    .B1(\__uuf__._0686_ ),
    .B2(\__uuf__._0687_ ),
    .X(\__uuf__._0691_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1641_ 
  (
    .A(\__uuf__._0664_ ),
    .B(\__uuf__._0688_ ),
    .C(\__uuf__._0691_ ),
    .X(\__uuf__._0692_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1642_ 
  (
    .A1(\__uuf__._0675_ ),
    .A2(\__uuf__._0688_ ),
    .B1(\__uuf__._0691_ ),
    .Y(\__uuf__._0693_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1643_ 
  (
    .A(\__uuf__._0682_ ),
    .B(\__uuf__._0692_ ),
    .C(\__uuf__._0693_ ),
    .X(\__uuf__._0016_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1644_ 
  (
    .A(\__uuf__._0014_ ),
    .Y(\__uuf__._0694_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1645_ 
  (
    .A(\__uuf__.multiplier.pp[8] ),
    .Y(\__uuf__._0695_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1646_ 
  (
    .A(\__uuf__._0514_ ),
    .X(\__uuf__._0696_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1647_ 
  (
    .A(\__BoundaryScanRegister_input_7__.dout ),
    .Y(\__uuf__._0697_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1648_ 
  (
    .A1(\__uuf__._0694_ ),
    .A2(\__uuf__._0695_ ),
    .B1(\__uuf__._0696_ ),
    .B2(\__uuf__._0697_ ),
    .X(\__uuf__._0698_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1649_ 
  (
    .A1(\__uuf__._0694_ ),
    .A2(\__uuf__._0695_ ),
    .B1(\__uuf__._0660_ ),
    .C1(\__uuf__._0698_ ),
    .X(\__uuf__._0699_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1650_ 
  (
    .A(\__uuf__._0699_ ),
    .Y(\__uuf__._0012_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1651_ 
  (
    .A1_N(\__uuf__._0694_ ),
    .A2_N(\__uuf__._0695_ ),
    .B1(\__uuf__._0694_ ),
    .B2(\__uuf__._0695_ ),
    .X(\__uuf__._0700_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1652_ 
  (
    .A(\__uuf__._0664_ ),
    .B(\__uuf__._0697_ ),
    .C(\__uuf__._0700_ ),
    .X(\__uuf__._0701_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1653_ 
  (
    .A1(\__uuf__._0675_ ),
    .A2(\__uuf__._0697_ ),
    .B1(\__uuf__._0700_ ),
    .Y(\__uuf__._0702_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1654_ 
  (
    .A(\__uuf__._0682_ ),
    .B(\__uuf__._0701_ ),
    .C(\__uuf__._0702_ ),
    .X(\__uuf__._0013_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1655_ 
  (
    .A(\__uuf__._0011_ ),
    .Y(\__uuf__._0703_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1656_ 
  (
    .A(\__uuf__.multiplier.pp[7] ),
    .Y(\__uuf__._0704_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1657_ 
  (
    .A(\__uuf__._0448_ ),
    .X(\__uuf__._0705_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1658_ 
  (
    .A(\__BoundaryScanRegister_input_6__.dout ),
    .Y(\__uuf__._0706_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1659_ 
  (
    .A1(\__uuf__._0703_ ),
    .A2(\__uuf__._0704_ ),
    .B1(\__uuf__._0696_ ),
    .B2(\__uuf__._0706_ ),
    .X(\__uuf__._0707_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1660_ 
  (
    .A1(\__uuf__._0703_ ),
    .A2(\__uuf__._0704_ ),
    .B1(\__uuf__._0705_ ),
    .C1(\__uuf__._0707_ ),
    .X(\__uuf__._0708_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1661_ 
  (
    .A(\__uuf__._0708_ ),
    .Y(\__uuf__._0009_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1662_ 
  (
    .A(\__uuf__._0487_ ),
    .X(\__uuf__._0709_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1663_ 
  (
    .A1_N(\__uuf__._0703_ ),
    .A2_N(\__uuf__._0704_ ),
    .B1(\__uuf__._0703_ ),
    .B2(\__uuf__._0704_ ),
    .X(\__uuf__._0710_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1664_ 
  (
    .A(\__uuf__._0709_ ),
    .B(\__uuf__._0706_ ),
    .C(\__uuf__._0710_ ),
    .X(\__uuf__._0711_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1665_ 
  (
    .A1(\__uuf__._0675_ ),
    .A2(\__uuf__._0706_ ),
    .B1(\__uuf__._0710_ ),
    .Y(\__uuf__._0712_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1666_ 
  (
    .A(\__uuf__._0682_ ),
    .B(\__uuf__._0711_ ),
    .C(\__uuf__._0712_ ),
    .X(\__uuf__._0010_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1667_ 
  (
    .A(\__uuf__._0008_ ),
    .Y(\__uuf__._0713_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1668_ 
  (
    .A(\__uuf__.multiplier.pp[6] ),
    .Y(\__uuf__._0714_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1669_ 
  (
    .A(\__BoundaryScanRegister_input_5__.dout ),
    .Y(\__uuf__._0715_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1670_ 
  (
    .A1(\__uuf__._0713_ ),
    .A2(\__uuf__._0714_ ),
    .B1(\__uuf__._0696_ ),
    .B2(\__uuf__._0715_ ),
    .X(\__uuf__._0716_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1671_ 
  (
    .A1(\__uuf__._0713_ ),
    .A2(\__uuf__._0714_ ),
    .B1(\__uuf__._0705_ ),
    .C1(\__uuf__._0716_ ),
    .X(\__uuf__._0717_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1672_ 
  (
    .A(\__uuf__._0717_ ),
    .Y(\__uuf__._0006_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1673_ 
  (
    .A1_N(\__uuf__._0713_ ),
    .A2_N(\__uuf__._0714_ ),
    .B1(\__uuf__._0713_ ),
    .B2(\__uuf__._0714_ ),
    .X(\__uuf__._0718_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1674_ 
  (
    .A(\__uuf__._0709_ ),
    .B(\__uuf__._0715_ ),
    .C(\__uuf__._0718_ ),
    .X(\__uuf__._0719_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1675_ 
  (
    .A(\__uuf__._0528_ ),
    .X(\__uuf__._0720_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1676_ 
  (
    .A1(\__uuf__._0720_ ),
    .A2(\__uuf__._0715_ ),
    .B1(\__uuf__._0718_ ),
    .Y(\__uuf__._0721_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1677_ 
  (
    .A(\__uuf__._0682_ ),
    .B(\__uuf__._0719_ ),
    .C(\__uuf__._0721_ ),
    .X(\__uuf__._0007_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1678_ 
  (
    .A(\__uuf__._0005_ ),
    .Y(\__uuf__._0722_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1679_ 
  (
    .A(\__uuf__.multiplier.pp[5] ),
    .Y(\__uuf__._0723_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1680_ 
  (
    .A(\__BoundaryScanRegister_input_4__.dout ),
    .Y(\__uuf__._0724_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1681_ 
  (
    .A1(\__uuf__._0722_ ),
    .A2(\__uuf__._0723_ ),
    .B1(\__uuf__._0696_ ),
    .B2(\__uuf__._0724_ ),
    .X(\__uuf__._0725_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1682_ 
  (
    .A1(\__uuf__._0722_ ),
    .A2(\__uuf__._0723_ ),
    .B1(\__uuf__._0705_ ),
    .C1(\__uuf__._0725_ ),
    .X(\__uuf__._0726_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1683_ 
  (
    .A(\__uuf__._0726_ ),
    .Y(\__uuf__._0003_ )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1684_ 
  (
    .A(\__uuf__._0807_ ),
    .X(\__uuf__._0727_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1685_ 
  (
    .A1_N(\__uuf__._0722_ ),
    .A2_N(\__uuf__._0723_ ),
    .B1(\__uuf__._0722_ ),
    .B2(\__uuf__._0723_ ),
    .X(\__uuf__._0728_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1686_ 
  (
    .A(\__uuf__._0709_ ),
    .B(\__uuf__._0724_ ),
    .C(\__uuf__._0728_ ),
    .X(\__uuf__._0729_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1687_ 
  (
    .A1(\__uuf__._0720_ ),
    .A2(\__uuf__._0724_ ),
    .B1(\__uuf__._0728_ ),
    .Y(\__uuf__._0730_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1688_ 
  (
    .A(\__uuf__._0727_ ),
    .B(\__uuf__._0729_ ),
    .C(\__uuf__._0730_ ),
    .X(\__uuf__._0004_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1689_ 
  (
    .A(\__uuf__._0002_ ),
    .Y(\__uuf__._0731_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1690_ 
  (
    .A(\__uuf__.multiplier.pp[4] ),
    .Y(\__uuf__._0732_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1691_ 
  (
    .A(\__BoundaryScanRegister_input_3__.dout ),
    .Y(\__uuf__._0733_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1692_ 
  (
    .A1(\__uuf__._0731_ ),
    .A2(\__uuf__._0732_ ),
    .B1(\__uuf__._0696_ ),
    .B2(\__uuf__._0733_ ),
    .X(\__uuf__._0734_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1693_ 
  (
    .A1(\__uuf__._0731_ ),
    .A2(\__uuf__._0732_ ),
    .B1(\__uuf__._0705_ ),
    .C1(\__uuf__._0734_ ),
    .X(\__uuf__._0735_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1694_ 
  (
    .A(\__uuf__._0735_ ),
    .Y(\__uuf__._0000_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1695_ 
  (
    .A1_N(\__uuf__._0731_ ),
    .A2_N(\__uuf__._0732_ ),
    .B1(\__uuf__._0731_ ),
    .B2(\__uuf__._0732_ ),
    .X(\__uuf__._0736_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1696_ 
  (
    .A(\__uuf__._0709_ ),
    .B(\__uuf__._0733_ ),
    .C(\__uuf__._0736_ ),
    .X(\__uuf__._0737_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1697_ 
  (
    .A1(\__uuf__._0720_ ),
    .A2(\__uuf__._0733_ ),
    .B1(\__uuf__._0736_ ),
    .Y(\__uuf__._0738_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1698_ 
  (
    .A(\__uuf__._0727_ ),
    .B(\__uuf__._0737_ ),
    .C(\__uuf__._0738_ ),
    .X(\__uuf__._0001_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1699_ 
  (
    .A(\__uuf__._0089_ ),
    .Y(\__uuf__._0739_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1700_ 
  (
    .A(\__uuf__.multiplier.pp[3] ),
    .Y(\__uuf__._0740_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1701_ 
  (
    .A(\__BoundaryScanRegister_input_2__.dout ),
    .Y(\__uuf__._0741_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1702_ 
  (
    .A1(\__uuf__._0739_ ),
    .A2(\__uuf__._0740_ ),
    .B1(\__uuf__._0491_ ),
    .B2(\__uuf__._0741_ ),
    .X(\__uuf__._0742_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1703_ 
  (
    .A1(\__uuf__._0739_ ),
    .A2(\__uuf__._0740_ ),
    .B1(\__uuf__._0705_ ),
    .C1(\__uuf__._0742_ ),
    .X(\__uuf__._0743_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1704_ 
  (
    .A(\__uuf__._0743_ ),
    .Y(\__uuf__._0087_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1705_ 
  (
    .A1_N(\__uuf__._0739_ ),
    .A2_N(\__uuf__._0740_ ),
    .B1(\__uuf__._0739_ ),
    .B2(\__uuf__._0740_ ),
    .X(\__uuf__._0744_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1706_ 
  (
    .A(\__uuf__._0709_ ),
    .B(\__uuf__._0741_ ),
    .C(\__uuf__._0744_ ),
    .X(\__uuf__._0745_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1707_ 
  (
    .A1(\__uuf__._0720_ ),
    .A2(\__uuf__._0741_ ),
    .B1(\__uuf__._0744_ ),
    .Y(\__uuf__._0746_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1708_ 
  (
    .A(\__uuf__._0727_ ),
    .B(\__uuf__._0745_ ),
    .C(\__uuf__._0746_ ),
    .X(\__uuf__._0088_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1709_ 
  (
    .A(\__uuf__._0086_ ),
    .Y(\__uuf__._0747_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1710_ 
  (
    .A(\__uuf__.multiplier.pp[2] ),
    .Y(\__uuf__._0748_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1711_ 
  (
    .A(\__BoundaryScanRegister_input_1__.dout ),
    .Y(\__uuf__._0749_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1712_ 
  (
    .A1(\__uuf__._0747_ ),
    .A2(\__uuf__._0748_ ),
    .B1(\__uuf__._0491_ ),
    .B2(\__uuf__._0749_ ),
    .X(\__uuf__._0750_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1713_ 
  (
    .A1(\__uuf__._0747_ ),
    .A2(\__uuf__._0748_ ),
    .B1(\__uuf__._0449_ ),
    .C1(\__uuf__._0750_ ),
    .X(\__uuf__._0751_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1714_ 
  (
    .A(\__uuf__._0751_ ),
    .Y(\__uuf__._0084_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1715_ 
  (
    .A1_N(\__uuf__._0747_ ),
    .A2_N(\__uuf__._0748_ ),
    .B1(\__uuf__._0747_ ),
    .B2(\__uuf__._0748_ ),
    .X(\__uuf__._0752_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1716_ 
  (
    .A(\__uuf__._0483_ ),
    .B(\__uuf__._0749_ ),
    .C(\__uuf__._0752_ ),
    .X(\__uuf__._0753_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1717_ 
  (
    .A1(\__uuf__._0720_ ),
    .A2(\__uuf__._0749_ ),
    .B1(\__uuf__._0752_ ),
    .Y(\__uuf__._0754_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1718_ 
  (
    .A(\__uuf__._0727_ ),
    .B(\__uuf__._0753_ ),
    .C(\__uuf__._0754_ ),
    .X(\__uuf__._0085_ )
  );


  sky130_fd_sc_hd__and2_4
  \__uuf__._1719_ 
  (
    .A(\__uuf__.multiplier.y ),
    .B(\__BoundaryScanRegister_input_31__.dout ),
    .X(\__uuf__._0755_ )
  );


  sky130_fd_sc_hd__o21a_4
  \__uuf__._1720_ 
  (
    .A1(\__uuf__.multiplier.tcmp.z ),
    .A2(\__uuf__._0755_ ),
    .B1(\__uuf__._0499_ ),
    .X(\__uuf__._0093_ )
  );


  sky130_fd_sc_hd__a21boi_4
  \__uuf__._1721_ 
  (
    .A1(\__uuf__.multiplier.tcmp.z ),
    .A2(\__uuf__._0755_ ),
    .B1_N(\__uuf__._0093_ ),
    .Y(\__uuf__._0092_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1722_ 
  (
    .A(\__uuf__.multiplier.csa0.sc ),
    .Y(\__uuf__._0756_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1723_ 
  (
    .A(\__uuf__.multiplier.csa0.y ),
    .Y(\__uuf__._0757_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1724_ 
  (
    .A(\__BoundaryScanRegister_input_0__.dout ),
    .Y(\__uuf__._0758_ )
  );


  sky130_fd_sc_hd__o22a_4
  \__uuf__._1725_ 
  (
    .A1(\__uuf__._0756_ ),
    .A2(\__uuf__._0757_ ),
    .B1(\__uuf__._0491_ ),
    .B2(\__uuf__._0758_ ),
    .X(\__uuf__._0759_ )
  );


  sky130_fd_sc_hd__a211o_4
  \__uuf__._1726_ 
  (
    .A1(\__uuf__._0756_ ),
    .A2(\__uuf__._0757_ ),
    .B1(\__uuf__._0449_ ),
    .C1(\__uuf__._0759_ ),
    .X(\__uuf__._0760_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1727_ 
  (
    .A(\__uuf__._0760_ ),
    .Y(\__uuf__._0090_ )
  );


  sky130_fd_sc_hd__a2bb2o_4
  \__uuf__._1728_ 
  (
    .A1_N(\__uuf__._0756_ ),
    .A2_N(\__uuf__._0757_ ),
    .B1(\__uuf__._0756_ ),
    .B2(\__uuf__._0757_ ),
    .X(\__uuf__._0761_ )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1729_ 
  (
    .A(\__uuf__._0483_ ),
    .B(\__uuf__._0758_ ),
    .C(\__uuf__._0761_ ),
    .X(\__uuf__._0762_ )
  );


  sky130_fd_sc_hd__o21ai_4
  \__uuf__._1730_ 
  (
    .A1(\__uuf__._0488_ ),
    .A2(\__uuf__._0758_ ),
    .B1(\__uuf__._0761_ ),
    .Y(\__uuf__._0763_ )
  );


  sky130_fd_sc_hd__and3_4
  \__uuf__._1731_ 
  (
    .A(\__uuf__._0727_ ),
    .B(\__uuf__._0762_ ),
    .C(\__uuf__._0763_ ),
    .X(\__uuf__._0091_ )
  );


  sky130_fd_sc_hd__and2_4
  \__uuf__._1732_ 
  (
    .A(\__BoundaryScanRegister_input_64__.dout ),
    .B(\__uuf__._0789_ ),
    .X(\__uuf__.fsm.newstate[0] )
  );


  sky130_fd_sc_hd__or3_4
  \__uuf__._1733_ 
  (
    .A(\__uuf__._0766_ ),
    .B(\__uuf__.fsm.state[1] ),
    .C(\__uuf__._0770_ ),
    .X(\__uuf__._0764_ )
  );


  sky130_fd_sc_hd__inv_2
  \__uuf__._1734_ 
  (
    .A(\__uuf__._0764_ ),
    .Y(\__uuf__._0765_ )
  );


  sky130_fd_sc_hd__o21a_4
  \__uuf__._1735_ 
  (
    .A1(done),
    .A2(\__uuf__._0765_ ),
    .B1(\__BoundaryScanRegister_input_64__.dout ),
    .X(\__uuf__.fsm.newstate[1] )
  );


  sky130_fd_sc_hd__buf_2
  \__uuf__._1736_ 
  (
    .A(\__uuf__._0794_ ),
    .X(\__uuf__._0360_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1737_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0342_),
    .Q(\__uuf__.shifter.shiftreg[0] ),
    .RESET_B(\__uuf__._0159_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1738_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0343_),
    .Q(\__uuf__.shifter.shiftreg[1] ),
    .RESET_B(\__uuf__._0160_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1739_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0344_),
    .Q(\__uuf__.shifter.shiftreg[2] ),
    .RESET_B(\__uuf__._0161_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1740_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0345_),
    .Q(\__uuf__.shifter.shiftreg[3] ),
    .RESET_B(\__uuf__._0162_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1741_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0346_),
    .Q(\__uuf__.shifter.shiftreg[4] ),
    .RESET_B(\__uuf__._0163_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1742_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0347_),
    .Q(\__uuf__.shifter.shiftreg[5] ),
    .RESET_B(\__uuf__._0164_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1743_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0348_),
    .Q(\__uuf__.shifter.shiftreg[6] ),
    .RESET_B(\__uuf__._0165_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1744_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0349_),
    .Q(\__uuf__.shifter.shiftreg[7] ),
    .RESET_B(\__uuf__._0166_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1745_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0350_),
    .Q(\__uuf__.shifter.shiftreg[8] ),
    .RESET_B(\__uuf__._0167_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1746_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0351_),
    .Q(\__uuf__.shifter.shiftreg[9] ),
    .RESET_B(\__uuf__._0168_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1747_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0352_),
    .Q(\__uuf__.shifter.shiftreg[10] ),
    .RESET_B(\__uuf__._0169_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1748_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0353_),
    .Q(\__uuf__.shifter.shiftreg[11] ),
    .RESET_B(\__uuf__._0170_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1749_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0354_),
    .Q(\__uuf__.shifter.shiftreg[12] ),
    .RESET_B(\__uuf__._0171_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1750_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0355_),
    .Q(\__uuf__.shifter.shiftreg[13] ),
    .RESET_B(\__uuf__._0172_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1751_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0356_),
    .Q(\__uuf__.shifter.shiftreg[14] ),
    .RESET_B(\__uuf__._0173_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1752_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0357_),
    .Q(\__uuf__.shifter.shiftreg[15] ),
    .RESET_B(\__uuf__._0174_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1753_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0358_),
    .Q(\__uuf__.shifter.shiftreg[16] ),
    .RESET_B(\__uuf__._0175_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1754_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0359_),
    .Q(\__uuf__.shifter.shiftreg[17] ),
    .RESET_B(\__uuf__._0176_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1755_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0360_),
    .Q(\__uuf__.shifter.shiftreg[18] ),
    .RESET_B(\__uuf__._0177_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1756_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0361_),
    .Q(\__uuf__.shifter.shiftreg[19] ),
    .RESET_B(\__uuf__._0178_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1757_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0362_),
    .Q(\__uuf__.shifter.shiftreg[20] ),
    .RESET_B(\__uuf__._0179_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1758_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0363_),
    .Q(\__uuf__.shifter.shiftreg[21] ),
    .RESET_B(\__uuf__._0180_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1759_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0364_),
    .Q(\__uuf__.shifter.shiftreg[22] ),
    .RESET_B(\__uuf__._0181_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1760_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0365_),
    .Q(\__uuf__.shifter.shiftreg[23] ),
    .RESET_B(\__uuf__._0182_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1761_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0366_),
    .Q(\__uuf__.shifter.shiftreg[24] ),
    .RESET_B(\__uuf__._0183_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1762_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0367_),
    .Q(\__uuf__.shifter.shiftreg[25] ),
    .RESET_B(\__uuf__._0184_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1763_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0368_),
    .Q(\__uuf__.shifter.shiftreg[26] ),
    .RESET_B(\__uuf__._0185_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1764_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0369_),
    .Q(\__uuf__.shifter.shiftreg[27] ),
    .RESET_B(\__uuf__._0186_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1765_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0370_),
    .Q(\__uuf__.shifter.shiftreg[28] ),
    .RESET_B(\__uuf__._0187_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1766_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0371_),
    .Q(\__uuf__.shifter.shiftreg[29] ),
    .RESET_B(\__uuf__._0188_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1767_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0372_),
    .Q(\__uuf__.shifter.shiftreg[30] ),
    .RESET_B(\__uuf__._0189_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1768_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0373_),
    .Q(\__uuf__.shifter.shiftreg[31] ),
    .RESET_B(\__uuf__._0190_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1769_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0374_),
    .Q(\__uuf__.shifter.shiftreg[32] ),
    .RESET_B(\__uuf__._0191_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1770_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0375_),
    .Q(\__uuf__.shifter.shiftreg[33] ),
    .RESET_B(\__uuf__._0192_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1771_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0376_),
    .Q(\__uuf__.shifter.shiftreg[34] ),
    .RESET_B(\__uuf__._0193_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1772_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0377_),
    .Q(\__uuf__.shifter.shiftreg[35] ),
    .RESET_B(\__uuf__._0194_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1773_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0378_),
    .Q(\__uuf__.shifter.shiftreg[36] ),
    .RESET_B(\__uuf__._0195_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1774_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0379_),
    .Q(\__uuf__.shifter.shiftreg[37] ),
    .RESET_B(\__uuf__._0196_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1775_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0380_),
    .Q(\__uuf__.shifter.shiftreg[38] ),
    .RESET_B(\__uuf__._0197_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1776_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0381_),
    .Q(\__uuf__.shifter.shiftreg[39] ),
    .RESET_B(\__uuf__._0198_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1777_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0382_),
    .Q(\__uuf__.shifter.shiftreg[40] ),
    .RESET_B(\__uuf__._0199_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1778_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0383_),
    .Q(\__uuf__.shifter.shiftreg[41] ),
    .RESET_B(\__uuf__._0200_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1779_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0384_),
    .Q(\__uuf__.shifter.shiftreg[42] ),
    .RESET_B(\__uuf__._0201_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1780_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0385_),
    .Q(\__uuf__.shifter.shiftreg[43] ),
    .RESET_B(\__uuf__._0202_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1781_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0386_),
    .Q(\__uuf__.shifter.shiftreg[44] ),
    .RESET_B(\__uuf__._0203_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1782_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0387_),
    .Q(\__uuf__.shifter.shiftreg[45] ),
    .RESET_B(\__uuf__._0204_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1783_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0388_),
    .Q(\__uuf__.shifter.shiftreg[46] ),
    .RESET_B(\__uuf__._0205_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1784_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0389_),
    .Q(\__uuf__.shifter.shiftreg[47] ),
    .RESET_B(\__uuf__._0206_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1785_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0390_),
    .Q(\__uuf__.shifter.shiftreg[48] ),
    .RESET_B(\__uuf__._0207_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1786_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0391_),
    .Q(\__uuf__.shifter.shiftreg[49] ),
    .RESET_B(\__uuf__._0208_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1787_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0392_),
    .Q(\__uuf__.shifter.shiftreg[50] ),
    .RESET_B(\__uuf__._0209_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1788_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0393_),
    .Q(\__uuf__.shifter.shiftreg[51] ),
    .RESET_B(\__uuf__._0210_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1789_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0394_),
    .Q(\__uuf__.shifter.shiftreg[52] ),
    .RESET_B(\__uuf__._0211_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1790_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0395_),
    .Q(\__uuf__.shifter.shiftreg[53] ),
    .RESET_B(\__uuf__._0212_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1791_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0396_),
    .Q(\__uuf__.shifter.shiftreg[54] ),
    .RESET_B(\__uuf__._0213_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1792_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0397_),
    .Q(\__uuf__.shifter.shiftreg[55] ),
    .RESET_B(\__uuf__._0214_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1793_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0398_),
    .Q(\__uuf__.shifter.shiftreg[56] ),
    .RESET_B(\__uuf__._0215_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1794_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0399_),
    .Q(\__uuf__.shifter.shiftreg[57] ),
    .RESET_B(\__uuf__._0216_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1795_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0400_),
    .Q(\__uuf__.shifter.shiftreg[58] ),
    .RESET_B(\__uuf__._0217_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1796_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0401_),
    .Q(\__uuf__.shifter.shiftreg[59] ),
    .RESET_B(\__uuf__._0218_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1797_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0402_),
    .Q(\__uuf__.shifter.shiftreg[60] ),
    .RESET_B(\__uuf__._0219_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1798_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0403_),
    .Q(\__uuf__.shifter.shiftreg[61] ),
    .RESET_B(\__uuf__._0220_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1799_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0404_),
    .Q(\__uuf__.shifter.shiftreg[62] ),
    .RESET_B(\__uuf__._0221_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1800_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0405_),
    .Q(\__uuf__.shifter.shiftreg[63] ),
    .RESET_B(\__uuf__._0222_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1801_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0406_),
    .Q(\__uuf__.multiplier.y ),
    .RESET_B(\__uuf__._0223_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1802_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0407_),
    .Q(\__uuf__.multiplier.pp[30] ),
    .RESET_B(\__uuf__._0224_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1803_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0408_),
    .Q(\__uuf__._0083_ ),
    .RESET_B(\__uuf__._0225_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1804_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0409_),
    .Q(\__uuf__.multiplier.pp[29] ),
    .RESET_B(\__uuf__._0226_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1805_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0410_),
    .Q(\__uuf__._0080_ ),
    .RESET_B(\__uuf__._0227_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1806_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0411_),
    .Q(\__uuf__.multiplier.pp[28] ),
    .RESET_B(\__uuf__._0228_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1807_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0412_),
    .Q(\__uuf__._0077_ ),
    .RESET_B(\__uuf__._0229_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1808_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0413_),
    .Q(\__uuf__.multiplier.pp[27] ),
    .RESET_B(\__uuf__._0230_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1809_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0414_),
    .Q(\__uuf__._0074_ ),
    .RESET_B(\__uuf__._0231_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1810_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0415_),
    .Q(\__uuf__.multiplier.pp[26] ),
    .RESET_B(\__uuf__._0232_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1811_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0416_),
    .Q(\__uuf__._0071_ ),
    .RESET_B(\__uuf__._0233_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1812_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0417_),
    .Q(\__uuf__.multiplier.pp[25] ),
    .RESET_B(\__uuf__._0234_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1813_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0418_),
    .Q(\__uuf__._0068_ ),
    .RESET_B(\__uuf__._0235_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1814_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0419_),
    .Q(\__uuf__.multiplier.pp[24] ),
    .RESET_B(\__uuf__._0236_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1815_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0420_),
    .Q(\__uuf__._0065_ ),
    .RESET_B(\__uuf__._0237_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1816_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0421_),
    .Q(\__uuf__.multiplier.pp[23] ),
    .RESET_B(\__uuf__._0238_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1817_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0422_),
    .Q(\__uuf__._0062_ ),
    .RESET_B(\__uuf__._0239_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1818_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0423_),
    .Q(\__uuf__.multiplier.pp[22] ),
    .RESET_B(\__uuf__._0240_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1819_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0424_),
    .Q(\__uuf__._0059_ ),
    .RESET_B(\__uuf__._0241_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1820_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0425_),
    .Q(\__uuf__.multiplier.pp[21] ),
    .RESET_B(\__uuf__._0242_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1821_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0426_),
    .Q(\__uuf__._0056_ ),
    .RESET_B(\__uuf__._0243_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1822_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0427_),
    .Q(\__uuf__.multiplier.pp[20] ),
    .RESET_B(\__uuf__._0244_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1823_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0428_),
    .Q(\__uuf__._0053_ ),
    .RESET_B(\__uuf__._0245_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1824_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0429_),
    .Q(\__uuf__.multiplier.pp[19] ),
    .RESET_B(\__uuf__._0246_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1825_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0430_),
    .Q(\__uuf__._0050_ ),
    .RESET_B(\__uuf__._0247_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1826_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0431_),
    .Q(\__uuf__.multiplier.pp[18] ),
    .RESET_B(\__uuf__._0248_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1827_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0432_),
    .Q(\__uuf__._0047_ ),
    .RESET_B(\__uuf__._0249_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1828_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0433_),
    .Q(\__uuf__.multiplier.pp[17] ),
    .RESET_B(\__uuf__._0250_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1829_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0434_),
    .Q(\__uuf__._0044_ ),
    .RESET_B(\__uuf__._0251_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1830_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0435_),
    .Q(\__uuf__.multiplier.pp[16] ),
    .RESET_B(\__uuf__._0252_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1831_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0436_),
    .Q(\__uuf__._0041_ ),
    .RESET_B(\__uuf__._0253_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1832_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0437_),
    .Q(\__uuf__.multiplier.pp[15] ),
    .RESET_B(\__uuf__._0254_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1833_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0438_),
    .Q(\__uuf__._0038_ ),
    .RESET_B(\__uuf__._0255_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1834_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0439_),
    .Q(\__uuf__.multiplier.pp[14] ),
    .RESET_B(\__uuf__._0256_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1835_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0440_),
    .Q(\__uuf__._0035_ ),
    .RESET_B(\__uuf__._0257_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1836_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0441_),
    .Q(\__uuf__.multiplier.pp[13] ),
    .RESET_B(\__uuf__._0258_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1837_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0442_),
    .Q(\__uuf__._0032_ ),
    .RESET_B(\__uuf__._0259_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1838_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0443_),
    .Q(\__uuf__.multiplier.pp[12] ),
    .RESET_B(\__uuf__._0260_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1839_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0444_),
    .Q(\__uuf__._0029_ ),
    .RESET_B(\__uuf__._0261_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1840_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0445_),
    .Q(\__uuf__.multiplier.pp[11] ),
    .RESET_B(\__uuf__._0262_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1841_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0446_),
    .Q(\__uuf__._0026_ ),
    .RESET_B(\__uuf__._0263_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1842_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0447_),
    .Q(\__uuf__.multiplier.pp[10] ),
    .RESET_B(\__uuf__._0264_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1843_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0448_),
    .Q(\__uuf__._0023_ ),
    .RESET_B(\__uuf__._0265_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1844_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0449_),
    .Q(\__uuf__.multiplier.pp[9] ),
    .RESET_B(\__uuf__._0266_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1845_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0450_),
    .Q(\__uuf__._0020_ ),
    .RESET_B(\__uuf__._0267_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1846_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0451_),
    .Q(\__uuf__.multiplier.pp[8] ),
    .RESET_B(\__uuf__._0268_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1847_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0452_),
    .Q(\__uuf__._0017_ ),
    .RESET_B(\__uuf__._0269_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1848_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0453_),
    .Q(\__uuf__.multiplier.pp[7] ),
    .RESET_B(\__uuf__._0270_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1849_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0454_),
    .Q(\__uuf__._0014_ ),
    .RESET_B(\__uuf__._0271_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1850_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0455_),
    .Q(\__uuf__.multiplier.pp[6] ),
    .RESET_B(\__uuf__._0272_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1851_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0456_),
    .Q(\__uuf__._0011_ ),
    .RESET_B(\__uuf__._0273_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1852_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0457_),
    .Q(\__uuf__.multiplier.pp[5] ),
    .RESET_B(\__uuf__._0274_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1853_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0458_),
    .Q(\__uuf__._0008_ ),
    .RESET_B(\__uuf__._0275_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1854_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0459_),
    .Q(\__uuf__.multiplier.pp[4] ),
    .RESET_B(\__uuf__._0276_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1855_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0460_),
    .Q(\__uuf__._0005_ ),
    .RESET_B(\__uuf__._0277_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1856_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0461_),
    .Q(\__uuf__.multiplier.pp[3] ),
    .RESET_B(\__uuf__._0278_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1857_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0260_),
    .Q(\__uuf__._0002_ ),
    .RESET_B(\__uuf__._0279_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1858_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0261_),
    .Q(\__uuf__.multiplier.pp[2] ),
    .RESET_B(\__uuf__._0280_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1859_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0262_),
    .Q(\__uuf__._0089_ ),
    .RESET_B(\__uuf__._0281_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1860_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0263_),
    .Q(\__uuf__.multiplier.csa0.y ),
    .RESET_B(\__uuf__._0282_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1861_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0264_),
    .Q(\__uuf__._0086_ ),
    .RESET_B(\__uuf__._0283_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1862_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0265_),
    .Q(\__uuf__.multiplier.pp[31] ),
    .RESET_B(\__uuf__._0284_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1863_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0266_),
    .Q(\__uuf__.multiplier.tcmp.z ),
    .RESET_B(\__uuf__._0285_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1864_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0267_),
    .Q(\__uuf__.multiplier.csa0.sum ),
    .RESET_B(\__uuf__._0286_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1865_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0268_),
    .Q(\__uuf__.multiplier.csa0.sc ),
    .RESET_B(\__uuf__._0287_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1866_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0269_),
    .Q(\__uuf__.fsm.state[0] ),
    .RESET_B(\__uuf__._0288_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1867_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0270_),
    .Q(\__uuf__.fsm.state[1] ),
    .RESET_B(\__uuf__._0289_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1868_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0271_),
    .Q(prod[0]),
    .RESET_B(\__uuf__._0290_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1869_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0272_),
    .Q(prod[1]),
    .RESET_B(\__uuf__._0291_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1870_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0273_),
    .Q(prod[2]),
    .RESET_B(\__uuf__._0292_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1871_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0274_),
    .Q(prod[3]),
    .RESET_B(\__uuf__._0293_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1872_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0275_),
    .Q(prod[4]),
    .RESET_B(\__uuf__._0294_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1873_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0276_),
    .Q(prod[5]),
    .RESET_B(\__uuf__._0295_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1874_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0277_),
    .Q(prod[6]),
    .RESET_B(\__uuf__._0296_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1875_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0278_),
    .Q(prod[7]),
    .RESET_B(\__uuf__._0297_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1876_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0279_),
    .Q(prod[8]),
    .RESET_B(\__uuf__._0298_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1877_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0280_),
    .Q(prod[9]),
    .RESET_B(\__uuf__._0299_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1878_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0281_),
    .Q(prod[10]),
    .RESET_B(\__uuf__._0300_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1879_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0282_),
    .Q(prod[11]),
    .RESET_B(\__uuf__._0301_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1880_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0283_),
    .Q(prod[12]),
    .RESET_B(\__uuf__._0302_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1881_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0284_),
    .Q(prod[13]),
    .RESET_B(\__uuf__._0303_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1882_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0285_),
    .Q(prod[14]),
    .RESET_B(\__uuf__._0304_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1883_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0286_),
    .Q(prod[15]),
    .RESET_B(\__uuf__._0305_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1884_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0287_),
    .Q(prod[16]),
    .RESET_B(\__uuf__._0306_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1885_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0288_),
    .Q(prod[17]),
    .RESET_B(\__uuf__._0307_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1886_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0289_),
    .Q(prod[18]),
    .RESET_B(\__uuf__._0308_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1887_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0290_),
    .Q(prod[19]),
    .RESET_B(\__uuf__._0309_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1888_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0291_),
    .Q(prod[20]),
    .RESET_B(\__uuf__._0310_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1889_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0292_),
    .Q(prod[21]),
    .RESET_B(\__uuf__._0311_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1890_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0293_),
    .Q(prod[22]),
    .RESET_B(\__uuf__._0312_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1891_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0294_),
    .Q(prod[23]),
    .RESET_B(\__uuf__._0313_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1892_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0295_),
    .Q(prod[24]),
    .RESET_B(\__uuf__._0314_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1893_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0296_),
    .Q(prod[25]),
    .RESET_B(\__uuf__._0315_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1894_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0297_),
    .Q(prod[26]),
    .RESET_B(\__uuf__._0316_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1895_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0298_),
    .Q(prod[27]),
    .RESET_B(\__uuf__._0317_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1896_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0299_),
    .Q(prod[28]),
    .RESET_B(\__uuf__._0318_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1897_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0300_),
    .Q(prod[29]),
    .RESET_B(\__uuf__._0319_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1898_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0301_),
    .Q(prod[30]),
    .RESET_B(\__uuf__._0320_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1899_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0302_),
    .Q(prod[31]),
    .RESET_B(\__uuf__._0321_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1900_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0303_),
    .Q(prod[32]),
    .RESET_B(\__uuf__._0322_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1901_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0304_),
    .Q(prod[33]),
    .RESET_B(\__uuf__._0323_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1902_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0305_),
    .Q(prod[34]),
    .RESET_B(\__uuf__._0324_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1903_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0306_),
    .Q(prod[35]),
    .RESET_B(\__uuf__._0325_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1904_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0307_),
    .Q(prod[36]),
    .RESET_B(\__uuf__._0326_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1905_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0308_),
    .Q(prod[37]),
    .RESET_B(\__uuf__._0327_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1906_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0309_),
    .Q(prod[38]),
    .RESET_B(\__uuf__._0328_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1907_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0310_),
    .Q(prod[39]),
    .RESET_B(\__uuf__._0329_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1908_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0311_),
    .Q(prod[40]),
    .RESET_B(\__uuf__._0330_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1909_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0312_),
    .Q(prod[41]),
    .RESET_B(\__uuf__._0331_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1910_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0313_),
    .Q(prod[42]),
    .RESET_B(\__uuf__._0332_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1911_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0314_),
    .Q(prod[43]),
    .RESET_B(\__uuf__._0333_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1912_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0315_),
    .Q(prod[44]),
    .RESET_B(\__uuf__._0334_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1913_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0316_),
    .Q(prod[45]),
    .RESET_B(\__uuf__._0335_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1914_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0317_),
    .Q(prod[46]),
    .RESET_B(\__uuf__._0336_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1915_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0318_),
    .Q(prod[47]),
    .RESET_B(\__uuf__._0337_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1916_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0319_),
    .Q(prod[48]),
    .RESET_B(\__uuf__._0338_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1917_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0320_),
    .Q(prod[49]),
    .RESET_B(\__uuf__._0339_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1918_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0321_),
    .Q(prod[50]),
    .RESET_B(\__uuf__._0340_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1919_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0322_),
    .Q(prod[51]),
    .RESET_B(\__uuf__._0341_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1920_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0323_),
    .Q(prod[52]),
    .RESET_B(\__uuf__._0342_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1921_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0324_),
    .Q(prod[53]),
    .RESET_B(\__uuf__._0343_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1922_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0325_),
    .Q(prod[54]),
    .RESET_B(\__uuf__._0344_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1923_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0326_),
    .Q(prod[55]),
    .RESET_B(\__uuf__._0345_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1924_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0327_),
    .Q(prod[56]),
    .RESET_B(\__uuf__._0346_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1925_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0328_),
    .Q(prod[57]),
    .RESET_B(\__uuf__._0347_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1926_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0329_),
    .Q(prod[58]),
    .RESET_B(\__uuf__._0348_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1927_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0330_),
    .Q(prod[59]),
    .RESET_B(\__uuf__._0349_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1928_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0331_),
    .Q(prod[60]),
    .RESET_B(\__uuf__._0350_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1929_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0332_),
    .Q(prod[61]),
    .RESET_B(\__uuf__._0351_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1930_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0333_),
    .Q(prod[62]),
    .RESET_B(\__uuf__._0352_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1931_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0334_),
    .Q(prod[63]),
    .RESET_B(\__uuf__._0353_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1932_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0335_),
    .Q(\__uuf__.count[0] ),
    .RESET_B(\__uuf__._0354_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1933_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0336_),
    .Q(\__uuf__.count[1] ),
    .RESET_B(\__uuf__._0355_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1934_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0337_),
    .Q(\__uuf__.count[2] ),
    .RESET_B(\__uuf__._0356_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1935_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0338_),
    .Q(\__uuf__.count[3] ),
    .RESET_B(\__uuf__._0357_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1936_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0339_),
    .Q(\__uuf__.count[4] ),
    .RESET_B(\__uuf__._0358_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1937_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0340_),
    .Q(\__uuf__.count[5] ),
    .RESET_B(\__uuf__._0359_ )
  );


  sky130_fd_sc_hd__dfrtp_4
  \__uuf__._1938_ 
  (
    .CLK(\__uuf__.__clk_source__ ),
    .D(_0341_),
    .Q(\__BoundaryScanRegister_output_65__.sin ),
    .RESET_B(\__uuf__._0360_ )
  );


endmodule



module tap_top
(
  tms_pad_i,
  tck_pad_i,
  trst_pad_i,
  tdi_pad_i,
  tdo_pad_o,
  tdo_padoe_o,
  shift_dr_o,
  pause_dr_o,
  update_dr_o,
  capture_dr_o,
  exit1_dr_o,
  exit2_dr_o,
  test_logic_reset_o,
  run_test_idle_o,
  extest_select_o,
  sample_preload_select_o,
  mbist_select_o,
  debug_select_o,
  preload_chain_o,
  tdo_o,
  debug_tdi_i,
  bs_chain_tdi_i,
  mbist_tdi_i,
  chain_tdi_i
);

  input tms_pad_i;
  input tck_pad_i;
  input trst_pad_i;
  input tdi_pad_i;
  output tdo_pad_o;
  output tdo_padoe_o;
  output shift_dr_o;
  output pause_dr_o;
  output update_dr_o;
  output capture_dr_o;
  output test_logic_reset_o;
  output run_test_idle_o;
  output exit1_dr_o;
  output exit2_dr_o;
  output extest_select_o;
  output sample_preload_select_o;
  output mbist_select_o;
  output debug_select_o;
  output preload_chain_o;
  output tdo_o;
  input debug_tdi_i;
  input bs_chain_tdi_i;
  input mbist_tdi_i;
  input chain_tdi_i;
  reg test_logic_reset;
  reg run_test_idle;
  reg select_dr_scan;
  reg capture_dr;
  reg shift_dr;
  reg exit1_dr;
  reg pause_dr;
  reg exit2_dr;
  reg update_dr;
  reg select_ir_scan;
  reg capture_ir;
  reg shift_ir;reg shift_ir_neg;
  reg exit1_ir;
  reg pause_ir;
  reg exit2_ir;
  reg update_ir;
  reg extest_select;
  reg sample_preload_select;
  reg idcode_select;
  reg mbist_select;
  reg debug_select;
  reg bypass_select;
  reg preload_chain_select;
  reg tdo_pad_o;
  reg tdo_padoe_o;
  reg tms_q1;reg tms_q2;reg tms_q3;reg tms_q4;
  wire tms_reset;
  assign tdo_o = tdi_pad_i;
  assign shift_dr_o = shift_dr;
  assign pause_dr_o = pause_dr;
  assign update_dr_o = update_dr;
  assign capture_dr_o = capture_dr;
  assign test_logic_reset_o = test_logic_reset;
  assign run_test_idle_o = run_test_idle;
  assign exit1_dr_o = exit1_dr;
  assign exit2_dr_o = exit2_dr;
  assign extest_select_o = extest_select;
  assign sample_preload_select_o = sample_preload_select;
  assign mbist_select_o = mbist_select;
  assign debug_select_o = debug_select;
  assign preload_chain_o = preload_chain_select;

  always @(posedge tck_pad_i) begin
    tms_q1 <= #1 tms_pad_i;
    tms_q2 <= #1 tms_q1;
    tms_q3 <= #1 tms_q2;
    tms_q4 <= #1 tms_q3;
  end

  assign tms_reset = tms_q1 & tms_q2 & tms_q3 & tms_q4 & tms_pad_i;

  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) test_logic_reset <= #1 1'b1; 
    else if(tms_reset) test_logic_reset <= #1 1'b1; 
    else begin
      if(tms_pad_i & (test_logic_reset | select_ir_scan)) test_logic_reset <= #1 1'b1; 
      else test_logic_reset <= #1 1'b0;
    end
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) run_test_idle <= #1 1'b0; 
    else if(tms_reset) run_test_idle <= #1 1'b0; 
    else if(~tms_pad_i & (test_logic_reset | run_test_idle | update_dr | update_ir)) run_test_idle <= #1 1'b1; 
    else run_test_idle <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) select_dr_scan <= #1 1'b0; 
    else if(tms_reset) select_dr_scan <= #1 1'b0; 
    else if(tms_pad_i & (run_test_idle | update_dr | update_ir)) select_dr_scan <= #1 1'b1; 
    else select_dr_scan <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) capture_dr <= #1 1'b0; 
    else if(tms_reset) capture_dr <= #1 1'b0; 
    else if(~tms_pad_i & select_dr_scan) capture_dr <= #1 1'b1; 
    else capture_dr <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) shift_dr <= #1 1'b0; 
    else if(tms_reset) shift_dr <= #1 1'b0; 
    else if(~tms_pad_i & (capture_dr | shift_dr | exit2_dr)) shift_dr <= #1 1'b1; 
    else shift_dr <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) exit1_dr <= #1 1'b0; 
    else if(tms_reset) exit1_dr <= #1 1'b0; 
    else if(tms_pad_i & (capture_dr | shift_dr)) exit1_dr <= #1 1'b1; 
    else exit1_dr <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) pause_dr <= #1 1'b0; 
    else if(tms_reset) pause_dr <= #1 1'b0; 
    else if(~tms_pad_i & (exit1_dr | pause_dr)) pause_dr <= #1 1'b1; 
    else pause_dr <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) exit2_dr <= #1 1'b0; 
    else if(tms_reset) exit2_dr <= #1 1'b0; 
    else if(tms_pad_i & pause_dr) exit2_dr <= #1 1'b1; 
    else exit2_dr <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) update_dr <= #1 1'b0; 
    else if(tms_reset) update_dr <= #1 1'b0; 
    else if(tms_pad_i & (exit1_dr | exit2_dr)) update_dr <= #1 1'b1; 
    else update_dr <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) select_ir_scan <= #1 1'b0; 
    else if(tms_reset) select_ir_scan <= #1 1'b0; 
    else if(tms_pad_i & select_dr_scan) select_ir_scan <= #1 1'b1; 
    else select_ir_scan <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) capture_ir <= #1 1'b0; 
    else if(tms_reset) capture_ir <= #1 1'b0; 
    else if(~tms_pad_i & select_ir_scan) capture_ir <= #1 1'b1; 
    else capture_ir <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) shift_ir <= #1 1'b0; 
    else if(tms_reset) shift_ir <= #1 1'b0; 
    else if(~tms_pad_i & (capture_ir | shift_ir | exit2_ir)) shift_ir <= #1 1'b1; 
    else shift_ir <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) exit1_ir <= #1 1'b0; 
    else if(tms_reset) exit1_ir <= #1 1'b0; 
    else if(tms_pad_i & (capture_ir | shift_ir)) exit1_ir <= #1 1'b1; 
    else exit1_ir <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) pause_ir <= #1 1'b0; 
    else if(tms_reset) pause_ir <= #1 1'b0; 
    else if(~tms_pad_i & (exit1_ir | pause_ir)) pause_ir <= #1 1'b1; 
    else pause_ir <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) exit2_ir <= #1 1'b0; 
    else if(tms_reset) exit2_ir <= #1 1'b0; 
    else if(tms_pad_i & pause_ir) exit2_ir <= #1 1'b1; 
    else exit2_ir <= #1 1'b0;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) update_ir <= #1 1'b0; 
    else if(tms_reset) update_ir <= #1 1'b0; 
    else if(tms_pad_i & (exit1_ir | exit2_ir)) update_ir <= #1 1'b1; 
    else update_ir <= #1 1'b0;
  end

  reg [4-1:0] jtag_ir;
  reg [4-1:0] latched_jtag_ir;reg [4-1:0] latched_jtag_ir_neg;
  reg instruction_tdo;

  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) jtag_ir[4-1:0] <= #1 4'b0; 
    else if(capture_ir) jtag_ir <= #1 4'b0101; 
    else if(shift_ir) jtag_ir[4-1:0] <= #1 { tdi_pad_i, jtag_ir[4-1:1] }; 
  end


  always @(negedge tck_pad_i) begin
    instruction_tdo <= #1 jtag_ir[0];
  end

  reg [31:0] idcode_reg;
  reg idcode_tdo;

  always @(posedge tck_pad_i) begin
    if(idcode_select & shift_dr) idcode_reg <= #1 { tdi_pad_i, idcode_reg[31:1] }; 
    else idcode_reg <= #1 32'h149511c3;
  end


  always @(negedge tck_pad_i) begin
    idcode_tdo <= #1 idcode_reg;
  end

  reg bypassed_tdo;
  reg bypass_reg;

  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) bypass_reg <= #1 1'b0; 
    else if(shift_dr) bypass_reg <= #1 tdi_pad_i; 
  end


  always @(negedge tck_pad_i) begin
    bypassed_tdo <= #1 bypass_reg;
  end


  always @(posedge tck_pad_i or posedge trst_pad_i) begin
    if(trst_pad_i) latched_jtag_ir <= #1 4'b0010; 
    else if(tms_reset) latched_jtag_ir <= #1 4'b0010; 
    else if(update_ir) latched_jtag_ir <= #1 jtag_ir; 
  end


  always @(latched_jtag_ir) begin
    extest_select = 1'b0;
    sample_preload_select = 1'b0;
    idcode_select = 1'b0;
    mbist_select = 1'b0;
    debug_select = 1'b0;
    bypass_select = 1'b0;
    preload_chain_select = 1'b0;
    case(latched_jtag_ir)
      4'b0000: extest_select = 1'b1;
      4'b0001: sample_preload_select = 1'b1;
      4'b0010: idcode_select = 1'b1;
      4'b1001: mbist_select = 1'b1;
      4'b1000: debug_select = 1'b1;
      4'b1111: bypass_select = 1'b1;
      4'b0011: preload_chain_select = 1'b1;
      default: bypass_select = 1'b1;
    endcase
  end


  always @(shift_ir_neg or exit1_ir or instruction_tdo or latched_jtag_ir_neg or idcode_tdo or debug_tdi_i or bs_chain_tdi_i or mbist_tdi_i or chain_tdi_i or bypassed_tdo) begin
    if(shift_ir_neg) tdo_pad_o = instruction_tdo; 
    else begin
      case(latched_jtag_ir_neg)
        4'b0010: tdo_pad_o = idcode_tdo;
        4'b1000: tdo_pad_o = debug_tdi_i;
        4'b0001: tdo_pad_o = bs_chain_tdi_i;
        4'b0000: tdo_pad_o = bs_chain_tdi_i;
        4'b1001: tdo_pad_o = mbist_tdi_i;
        4'b0011: tdo_pad_o = chain_tdi_i;
        default: tdo_pad_o = bypassed_tdo;
      endcase
    end
  end


  always @(negedge tck_pad_i) begin
    tdo_padoe_o <= #1 shift_ir | shift_dr | pause_dr & debug_select;
  end


  always @(negedge tck_pad_i) begin
    shift_ir_neg <= #1 shift_ir;
    latched_jtag_ir_neg <= #1 latched_jtag_ir;
  end


endmodule

module spm_top
(
  mc,
  mp,
  clk,
  rst,
  prod,
  start,
  done,
  tms,
  tck,
  tdi,
  tdo,
  trst,
  tdo_paden_o
);

  input tms;
  input tck;
  input tdi;
  output tdo;
  output tdo_paden_o;
  input trst;
  input [31:0] mc;
  input [31:0] mp;
  input clk;
  input rst;
  input start;
  output [63:0] prod;
  output done;
  wire tdo_pad_o;
  wire tdo_paden_o;
  wire tms;
  wire tdi;
  wire trst;
  wire sin;
  wire sout;
  wire shift;
  wire test;

  tap_wrapper
  __tap_wrapper__
  (
    .tms(tms),
    .tck(tck),
    .trst(trst),
    .tdi(tdi),
    .tdo_pad_o(tdo),
    .tdo_paden_o(tdo_paden_o),
    .sin(sin),
    .sout(sout),
    .test(test),
    .shift(shift)
  );


  __DESIGN__UNDER__TEST__
  __dut__
  (
    .mc(mc),
    .mp(mp),
    .clk(clk),
    .rst(rst),
    .start(start),
    .sin(sin),
    .shift(shift),
    .tck(tck),
    .test(test),
    .prod(prod),
    .done(done),
    .sout(sout)
  );


endmodule


