* NGSPICE file created from spm_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt spm_top clk done mc[0] mc[10] mc[11] mc[12] mc[13] mc[14] mc[15] mc[16] mc[17]
+ mc[18] mc[19] mc[1] mc[20] mc[21] mc[22] mc[23] mc[24] mc[25] mc[26] mc[27] mc[28]
+ mc[29] mc[2] mc[30] mc[31] mc[3] mc[4] mc[5] mc[6] mc[7] mc[8] mc[9] mp[0] mp[10]
+ mp[11] mp[12] mp[13] mp[14] mp[15] mp[16] mp[17] mp[18] mp[19] mp[1] mp[20] mp[21]
+ mp[22] mp[23] mp[24] mp[25] mp[26] mp[27] mp[28] mp[29] mp[2] mp[30] mp[31] mp[3]
+ mp[4] mp[5] mp[6] mp[7] mp[8] mp[9] prod[0] prod[10] prod[11] prod[12] prod[13]
+ prod[14] prod[15] prod[16] prod[17] prod[18] prod[19] prod[1] prod[20] prod[21]
+ prod[22] prod[23] prod[24] prod[25] prod[26] prod[27] prod[28] prod[29] prod[2]
+ prod[30] prod[31] prod[32] prod[33] prod[34] prod[35] prod[36] prod[37] prod[38]
+ prod[39] prod[3] prod[40] prod[41] prod[42] prod[43] prod[44] prod[45] prod[46]
+ prod[47] prod[48] prod[49] prod[4] prod[50] prod[51] prod[52] prod[53] prod[54]
+ prod[55] prod[56] prod[57] prod[58] prod[59] prod[5] prod[60] prod[61] prod[62]
+ prod[63] prod[6] prod[7] prod[8] prod[9] rst start tck tdi tdo tdo_paden_o tms trst
+ VPWR VGND
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1505__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1240__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1506_ __dut__._1709_/X __dut__.__uuf__._1494_/X __dut__._1174_/B
+ __dut__.__uuf__._1495_/X VGND VGND VPWR VPWR __dut__.__uuf__._1506_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1437_ __dut__.__uuf__._1483_/A VGND VGND VPWR VPWR __dut__.__uuf__._1437_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1622_ __dut__._1766_/A __dut__._1808_/Q VGND VGND VPWR VPWR __dut__._1622_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1368_ __dut__._1232_/B VGND VGND VPWR VPWR __dut__.__uuf__._1368_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_14_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2200_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1299_ __dut__.__uuf__._1324_/A VGND VGND VPWR VPWR __dut__.__uuf__._1299_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1553_ __dut__._1543_/Y mc[11] __dut__._1552_/X VGND VGND VPWR VPWR __dut__._1553_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1484_ rst VGND VGND VPWR VPWR __dut__._1484_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1415__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1047__A __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_294_ _313_/CLK _294_/D trst VGND VGND VPWR VPWR _294_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__290__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__.__uuf__._2202__CLK __dut__.__uuf__._2210_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1222_ __dut__.__uuf__._1233_/A VGND VGND VPWR VPWR __dut__.__uuf__._1222_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1153_ __dut__.__uuf__._1212_/A VGND VGND VPWR VPWR __dut__.__uuf__._1153_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1084_ __dut__.__uuf__._1084_/A VGND VGND VPWR VPWR __dut__.__uuf__._1084_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_70_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1986_ __dut__.__uuf__._1986_/A VGND VGND VPWR VPWR __dut__._1125_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0984_ __dut__._0984_/A __dut__._1908_/Q VGND VGND VPWR VPWR __dut__._0984_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1605_ __dut__._1543_/Y mc[23] __dut__._1604_/X VGND VGND VPWR VPWR __dut__._1605_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1536_ rst VGND VGND VPWR VPWR __dut__._1536_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1467_ rst VGND VGND VPWR VPWR __dut__._1467_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1398_ __dut__._1408_/A __dut__._1398_/B VGND VGND VPWR VPWR __dut__._1398_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_61_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_12_0_tck clkbuf_3_6_0_tck/X VGND VGND VPWR VPWR __dut__._1902_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1837__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_277_ _313_/CLK _277_/D VGND VGND VPWR VPWR _277_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_156_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._0894__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1840_ __dut__.__uuf__._1883_/A __dut__.__uuf__._1840_/B __dut__.__uuf__._1840_/C
+ VGND VGND VPWR VPWR __dut__._1067_/A2 sky130_fd_sc_hd__and3_4
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1771_ __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR __dut__.__uuf__._1771_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._2185_ __dut__.__uuf__._2194_/CLK __dut__._1359_/X __dut__.__uuf__._1130_/X
+ VGND VGND VPWR VPWR prod[45] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1205_ __dut__.__uuf__._1249_/A VGND VGND VPWR VPWR __dut__.__uuf__._1205_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1143__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1136_ __dut__.__uuf__._1124_/X __dut__.__uuf__._1135_/X prod[44]
+ prod[45] __dut__.__uuf__._1131_/X VGND VGND VPWR VPWR __dut__._1357_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1067_ __dut__.__uuf__._2008_/A VGND VGND VPWR VPWR __dut__.__uuf__._1084_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1321_ __dut__._1339_/A1 __dut__._1321_/A2 __dut__._1320_/X VGND VGND VPWR
+ VPWR __dut__._1321_/X sky130_fd_sc_hd__a21o_4
X__dut__._1252_ __dut__._1408_/A __dut__._1252_/B VGND VGND VPWR VPWR __dut__._1252_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1183_ __dut__._1187_/A1 __dut__._1183_/A2 __dut__._1182_/X VGND VGND VPWR
+ VPWR __dut__._1183_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1969_ __dut__.__uuf__._1936_/X __dut__.__uuf__._1968_/B __dut__.__uuf__._1968_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1970_/C sky130_fd_sc_hd__o21ai_4
X_200_ _203_/A VGND VGND VPWR VPWR _200_/X sky130_fd_sc_hd__buf_2
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_131_ _309_/Q VGND VGND VPWR VPWR _131_/Y sky130_fd_sc_hd__inv_2
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_1_0_tck clkbuf_3_1_0_tck/A VGND VGND VPWR VPWR clkbuf_4_3_0_tck/A sky130_fd_sc_hd__clkbuf_1
Xpsn_inst_psn_buff_90 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1405_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._0967_ __dut__._0967_/A1 prod[15] __dut__._0966_/X VGND VGND VPWR VPWR __dut__._1900_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0898_ __dut__._1378_/A __dut__._1865_/Q VGND VGND VPWR VPWR __dut__._0898_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1685__A2 mp[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1519_ rst VGND VGND VPWR VPWR __dut__._1519_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1373__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1125__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1513__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1823_ __dut__.__uuf__._1823_/A VGND VGND VPWR VPWR __dut__._1065_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1754_ __dut__._1601_/X VGND VGND VPWR VPWR __dut__.__uuf__._1760_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1685_ __dut__.__uuf__._1685_/A VGND VGND VPWR VPWR __dut__.__uuf__._1923_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1870_ __dut__._1915_/CLK __dut__._1870_/D __dut__._1459_/Y VGND VGND VPWR
+ VPWR __dut__._1870_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2070__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2168_ __dut__.__uuf__._2169_/CLK __dut__._1325_/X __dut__.__uuf__._1182_/X
+ VGND VGND VPWR VPWR prod[28] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1119_ __dut__.__uuf__._1162_/A VGND VGND VPWR VPWR __dut__.__uuf__._1130_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2099_ __dut__.__uuf__._2164_/CLK __dut__._1187_/X __dut__.__uuf__._1470_/X
+ VGND VGND VPWR VPWR __dut__._1188_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1304_ __dut__._1304_/A prod[17] VGND VGND VPWR VPWR __dut__._1304_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1423__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_57_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1235_ __dut__._1787_/A1 __dut__._1235_/A2 __dut__._1234_/X VGND VGND VPWR
+ VPWR __dut__._1235_/X sky130_fd_sc_hd__a21o_4
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1166_ __dut__._1766_/A __dut__._1166_/B VGND VGND VPWR VPWR __dut__._1166_/X
+ sky130_fd_sc_hd__and2_4
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1097_ __dut__._1129_/A1 __dut__._1097_/A2 __dut__._1096_/X VGND VGND VPWR
+ VPWR __dut__._1097_/X sky130_fd_sc_hd__a21o_4
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1355__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1107__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_119_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2093__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1470_ __dut__.__uuf__._1486_/A VGND VGND VPWR VPWR __dut__.__uuf__._1470_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1508__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2022_ __dut__.__uuf__._2049_/CLK __dut__._1033_/X __dut__.__uuf__._1640_/X
+ VGND VGND VPWR VPWR __dut__._1034_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1649__A2 mp[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1020_ __dut__._1128_/A __dut__._1020_/B VGND VGND VPWR VPWR __dut__._1020_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_52_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1806_ __dut__.__uuf__._1828_/A __dut__.__uuf__._1806_/B __dut__.__uuf__._1806_/C
+ VGND VGND VPWR VPWR __dut__._1055_/A2 sky130_fd_sc_hd__and3_4
XANTENNA___dut__._1585__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1737_ __dut__.__uuf__._1731_/Y __dut__.__uuf__._1732_/Y __dut__.__uuf__._1731_/Y
+ __dut__.__uuf__._1732_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1738_/C sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1668_ __dut__.__uuf__._1868_/A VGND VGND VPWR VPWR __dut__.__uuf__._1692_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1853_ clkbuf_4_5_0_tck/X __dut__._1853_/D __dut__._1476_/Y VGND VGND VPWR
+ VPWR __dut__._1853_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1599_ __dut__.__uuf__._1599_/A VGND VGND VPWR VPWR __dut__.__uuf__._1599_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1418__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1784_ __dut__._1788_/A __dut__._1850_/Q VGND VGND VPWR VPWR __dut__._1784_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_0_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1218_ __dut__._1786_/A __dut__._1218_/B VGND VGND VPWR VPWR __dut__._1218_/X
+ sky130_fd_sc_hd__and2_4
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1149_ __dut__._1151_/A1 __dut__._1149_/A2 __dut__._1148_/X VGND VGND VPWR
+ VPWR __dut__._1149_/X sky130_fd_sc_hd__a21o_4
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1328__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1567__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1522_ __dut__.__uuf__._1529_/A VGND VGND VPWR VPWR __dut__.__uuf__._1522_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1453_ __dut__._1769_/X __dut__.__uuf__._1451_/X __dut__._1200_/B
+ __dut__.__uuf__._1452_/X VGND VGND VPWR VPWR __dut__.__uuf__._1453_/X sky130_fd_sc_hd__o22a_4
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1384_ __dut__.__uuf__._1393_/A VGND VGND VPWR VPWR __dut__.__uuf__._1384_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1238__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2005_ __dut__.__uuf__._2005_/A __dut__._1138_/B __dut__.__uuf__._2005_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2006_/A sky130_fd_sc_hd__or3_4
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1003_ __dut__._1339_/A1 prod[33] __dut__._1002_/X VGND VGND VPWR VPWR __dut__._1918_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1870__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1905_ clkbuf_4_9_0_tck/X __dut__._1905_/D __dut__._1424_/Y VGND VGND VPWR
+ VPWR __dut__._1905_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1836_ __dut__._1902_/CLK __dut__._1836_/D __dut__._1493_/Y VGND VGND VPWR
+ VPWR __dut__._1836_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1767_ __dut__._1767_/A1 __dut__._1765_/X __dut__._1766_/X VGND VGND VPWR
+ VPWR __dut__._1845_/D sky130_fd_sc_hd__a21o_4
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1698_ __dut__._1766_/A __dut__._1827_/Q VGND VGND VPWR VPWR __dut__._1698_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_48_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__127__A tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1549__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1081__B2 __dut__.__uuf__._1069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1058__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1721__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1521__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1893__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1505_ __dut__.__uuf__._1566_/A VGND VGND VPWR VPWR __dut__.__uuf__._1505_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1436_ __dut__.__uuf__._1442_/A VGND VGND VPWR VPWR __dut__.__uuf__._1436_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1621_ __dut__._1543_/Y mc[27] __dut__._1620_/X VGND VGND VPWR VPWR __dut__._1621_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1367_ __dut__.__uuf__._1367_/A VGND VGND VPWR VPWR __dut__.__uuf__._1367_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1552_ __dut__._1788_/A __dut__._1792_/Q VGND VGND VPWR VPWR __dut__._1552_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1298_ __dut__.__uuf__._1401_/A VGND VGND VPWR VPWR __dut__.__uuf__._1324_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0___dut__.__uuf__.__clk_source__/X sky130_fd_sc_hd__clkbuf_1
X__dut__._1483_ rst VGND VGND VPWR VPWR __dut__._1483_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1431__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_293_ _306_/CLK _293_/D trst VGND VGND VPWR VPWR _293_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1819_ clkbuf_4_6_0_tck/X __dut__._1819_/D __dut__._1510_/Y VGND VGND VPWR
+ VPWR __dut__._1819_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1606__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1238__A __dut__.__uuf__._1450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_101_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._1221_ __dut__.__uuf__._1236_/A VGND VGND VPWR VPWR __dut__.__uuf__._1233_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_101_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1152_ __dut__.__uuf__._1226_/A VGND VGND VPWR VPWR __dut__.__uuf__._1212_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_101_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1083_ __dut__.__uuf__._1075_/X __dut__.__uuf__._2003_/A prod[61]
+ prod[62] __dut__.__uuf__._1069_/X VGND VGND VPWR VPWR __dut__._1391_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1516__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1985_ __dut__.__uuf__._1981_/Y __dut__.__uuf__._1982_/Y __dut__.__uuf__._1941_/X
+ __dut__.__uuf__._1984_/X VGND VGND VPWR VPWR __dut__.__uuf__._1986_/A sky130_fd_sc_hd__a211o_4
XFILLER_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__308__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0983_ __dut__._0983_/A1 prod[23] __dut__._0982_/X VGND VGND VPWR VPWR __dut__._1908_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1419_ __dut__._1212_/B VGND VGND VPWR VPWR __dut__.__uuf__._1419_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1604_ __dut__._1788_/A __dut__._1805_/Q VGND VGND VPWR VPWR __dut__._1604_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1535_ rst VGND VGND VPWR VPWR __dut__._1535_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1426__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1466_ rst VGND VGND VPWR VPWR __dut__._1466_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1397_ __dut__._1409_/A1 __dut__._1397_/A2 __dut__._1396_/X VGND VGND VPWR
+ VPWR __dut__._1397_/X sky130_fd_sc_hd__a21o_4
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_276_ _314_/CLK _276_/D VGND VGND VPWR VPWR _276_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1336__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_149_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1770_ __dut__.__uuf__._1804_/A __dut__.__uuf__._1770_/B __dut__.__uuf__._1770_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1773_/B sky130_fd_sc_hd__or3_4
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2184_ __dut__.__uuf__._2194_/CLK __dut__._1357_/X __dut__.__uuf__._1134_/X
+ VGND VGND VPWR VPWR prod[44] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1204_ __dut__.__uuf__._1204_/A VGND VGND VPWR VPWR __dut__.__uuf__._1204_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1135_ __dut__.__uuf__._1149_/A VGND VGND VPWR VPWR __dut__.__uuf__._1135_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1320_ __dut__._1378_/A prod[25] VGND VGND VPWR VPWR __dut__._1320_/X sky130_fd_sc_hd__and2_4
XFILLER_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1066_ __dut__.__uuf__._1061_/B __dut__.__uuf__._1064_/X __dut__.__uuf__._1054_/X
+ __dut__._1400_/B __dut__.__uuf__._1314_/A VGND VGND VPWR VPWR __dut__._1399_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1251_ __dut__._1787_/A1 __dut__._1251_/A2 __dut__._1250_/X VGND VGND VPWR
+ VPWR __dut__._1251_/X sky130_fd_sc_hd__a21o_4
X__dut__._1182_ __dut__._1770_/A __dut__._1182_/B VGND VGND VPWR VPWR __dut__._1182_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1968_ __dut__.__uuf__._1968_/A __dut__.__uuf__._1968_/B __dut__.__uuf__._1968_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1970_/B sky130_fd_sc_hd__or3_4
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1899_ __dut__.__uuf__._1896_/Y __dut__.__uuf__._1897_/Y __dut__.__uuf__._1853_/X
+ __dut__.__uuf__._1903_/B VGND VGND VPWR VPWR __dut__.__uuf__._1899_/X sky130_fd_sc_hd__o22a_4
X_130_ _130_/A VGND VGND VPWR VPWR _314_/D sky130_fd_sc_hd__inv_2
XFILLER_7_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__280__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_91 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1409_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._0966_ __dut__._1324_/A __dut__._1899_/Q VGND VGND VPWR VPWR __dut__._0966_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_80 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1151_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._0897_ __dut__._1383_/A1 prod[45] __dut__._0896_/X VGND VGND VPWR VPWR __dut__._1865_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_78_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1156__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._0893__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1518_ rst VGND VGND VPWR VPWR __dut__._1518_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1449_ rst VGND VGND VPWR VPWR __dut__._1449_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1804__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1516__A __dut__.__uuf__._1720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_259_ _194_/A _259_/D VGND VGND VPWR VPWR _259_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__.__uuf__._1251__A __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1822_ __dut__.__uuf__._1818_/Y __dut__.__uuf__._1819_/Y __dut__.__uuf__._1776_/X
+ __dut__.__uuf__._1821_/X VGND VGND VPWR VPWR __dut__.__uuf__._1823_/A sky130_fd_sc_hd__a211o_4
XFILLER_40_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1753_ __dut__._1036_/B VGND VGND VPWR VPWR __dut__.__uuf__._1753_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._0939__A2 prod[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1684_ __dut__._1012_/B VGND VGND VPWR VPWR __dut__.__uuf__._1684_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_11_0_tck clkbuf_3_5_0_tck/X VGND VGND VPWR VPWR __dut__._1919_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_87_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2167_ __dut__.__uuf__._2169_/CLK __dut__._1323_/X __dut__.__uuf__._1185_/X
+ VGND VGND VPWR VPWR prod[27] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._0875__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1118_ __dut__.__uuf__._1109_/X __dut__.__uuf__._1106_/X prod[50]
+ prod[51] __dut__.__uuf__._1117_/X VGND VGND VPWR VPWR __dut__._1369_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2098_ __dut__.__uuf__._2164_/CLK __dut__._1185_/X __dut__.__uuf__._1476_/X
+ VGND VGND VPWR VPWR __dut__._1186_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1049_ __dut__._1408_/B __dut__.__uuf__._1052_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1049_/X sky130_fd_sc_hd__or2_4
X__dut__._1303_ __dut__._1319_/A1 __dut__._1303_/A2 __dut__._1302_/X VGND VGND VPWR
+ VPWR __dut__._1303_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1704__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1234_ __dut__._1786_/A __dut__._1234_/B VGND VGND VPWR VPWR __dut__._1234_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1165_ __dut__._1165_/A1 __dut__._1165_/A2 __dut__._1164_/X VGND VGND VPWR
+ VPWR __dut__._1165_/X sky130_fd_sc_hd__a21o_4
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1096_ __dut__._1678_/A __dut__._1096_/B VGND VGND VPWR VPWR __dut__._1096_/X
+ sky130_fd_sc_hd__and2_4
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._0949_ __dut__._0949_/A1 prod[6] __dut__._0948_/X VGND VGND VPWR VPWR __dut__._1891_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1614__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1043__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2021_ __dut__.__uuf__._2049_/CLK __dut__._1031_/X __dut__.__uuf__._1641_/X
+ VGND VGND VPWR VPWR __dut__._1032_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1524__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_tck clkbuf_3_1_0_tck/A VGND VGND VPWR VPWR clkbuf_4_1_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1805_ __dut__.__uuf__._1771_/X __dut__.__uuf__._1804_/B __dut__.__uuf__._1804_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1806_/C sky130_fd_sc_hd__o21ai_4
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1736_ __dut__.__uuf__._1736_/A VGND VGND VPWR VPWR __dut__._1033_/A2
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1585__A2 mc[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1667_ __dut__.__uuf__._1908_/A VGND VGND VPWR VPWR __dut__.__uuf__._1868_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1598_ __dut__.__uuf__._1599_/A VGND VGND VPWR VPWR __dut__.__uuf__._1598_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1852_ __dut__._1410_/B __dut__._1852_/D __dut__._1477_/Y VGND VGND VPWR
+ VPWR __dut__._1852_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1783_ __dut__._1787_/A1 __dut__._1781_/X __dut__._1782_/X VGND VGND VPWR
+ VPWR __dut__._1849_/D sky130_fd_sc_hd__a21o_4
XFILLER_0_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1434__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1217_ __dut__._1787_/A1 __dut__._1217_/A2 __dut__._1216_/X VGND VGND VPWR
+ VPWR __dut__._1217_/X sky130_fd_sc_hd__a21o_4
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1025__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1148_ __dut__._1150_/A __dut__._1148_/B VGND VGND VPWR VPWR __dut__._1148_/X
+ sky130_fd_sc_hd__and2_4
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1079_ __dut__._1129_/A1 __dut__._1079_/A2 __dut__._1078_/X VGND VGND VPWR
+ VPWR __dut__._1079_/X sky130_fd_sc_hd__a21o_4
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_131_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1521_ __dut__.__uuf__._1509_/X __dut__.__uuf__._1505_/X __dut__._1166_/B
+ __dut__.__uuf__._1514_/X __dut__.__uuf__._1520_/X VGND VGND VPWR VPWR __dut__._1165_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1452_ __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR __dut__.__uuf__._1452_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1519__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1383_ __dut__.__uuf__._1380_/X __dut__.__uuf__._1382_/X __dut__._1226_/B
+ __dut__.__uuf__._1380_/X VGND VGND VPWR VPWR __dut__._1225_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._2004_ __dut__._1785_/X __dut__.__uuf__._2004_/B VGND VGND VPWR VPWR
+ __dut__._1135_/A2 sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1254__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1255__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1002_ __dut__._1002_/A __dut__._1917_/Q VGND VGND VPWR VPWR __dut__._1002_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1007__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1719_ __dut__._1024_/B VGND VGND VPWR VPWR __dut__.__uuf__._1719_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1904_ clkbuf_4_9_0_tck/X __dut__._1904_/D __dut__._1425_/Y VGND VGND VPWR
+ VPWR __dut__._1904_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1429__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1835_ __dut__._1902_/CLK __dut__._1835_/D __dut__._1494_/Y VGND VGND VPWR
+ VPWR __dut__._1835_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1766_ __dut__._1766_/A __dut__._1834_/Q VGND VGND VPWR VPWR __dut__._1766_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1697_ __dut__._1543_/Y mp[12] __dut__._1696_/X VGND VGND VPWR VPWR __dut__._1697_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_48_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_3_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1164__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2083__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1549__A2 mc[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1081__A2 __dut__.__uuf__._2003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1721__A2 mc[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1237__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1504_ __dut__.__uuf__._1508_/A VGND VGND VPWR VPWR __dut__.__uuf__._1504_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1435_ __dut__.__uuf__._1070_/X __dut__.__uuf__._1434_/X __dut__._1204_/B
+ __dut__.__uuf__._1070_/X VGND VGND VPWR VPWR __dut__._1203_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1620_ __dut__._1788_/A __dut__._1809_/Q VGND VGND VPWR VPWR __dut__._1620_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1366_ __dut__.__uuf__._1354_/X __dut__.__uuf__._1364_/X __dut__._1232_/B
+ __dut__.__uuf__._1365_/X VGND VGND VPWR VPWR __dut__._1231_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1551_ __dut__._1767_/A1 __dut__._1549_/X __dut__._1550_/X VGND VGND VPWR
+ VPWR __dut__._1791_/D sky130_fd_sc_hd__a21o_4
XANTENNA_clkbuf_0___dut__.__uuf__.__clk_source___A __dut__._1411_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1297_ __dut__.__uuf__._1400_/A VGND VGND VPWR VPWR __dut__.__uuf__._1297_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_85_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1482_ rst VGND VGND VPWR VPWR __dut__._1482_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1712__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_292_ _306_/CLK _292_/D trst VGND VGND VPWR VPWR _292_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_psn_inst_psn_buff_32_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1818_ clkbuf_4_7_0_tck/X __dut__._1818_/D __dut__._1511_/Y VGND VGND VPWR
+ VPWR __dut__._1818_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._0998__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1749_ __dut__._1543_/Y mp[24] __dut__._1748_/X VGND VGND VPWR VPWR __dut__._1749_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1219__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1622__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1220_ __dut__.__uuf__._1212_/X __dut__.__uuf__._1209_/X prod[15]
+ prod[16] __dut__.__uuf__._1219_/X VGND VGND VPWR VPWR __dut__._1299_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1151_ __dut__.__uuf__._1159_/A VGND VGND VPWR VPWR __dut__.__uuf__._1151_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1082_ __dut__.__uuf__._1084_/A VGND VGND VPWR VPWR __dut__.__uuf__._1082_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_67_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1860__CLK __dut__._1917_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1532__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1164__A __dut__.__uuf__._1450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1984_ __dut__.__uuf__._1981_/Y __dut__.__uuf__._1982_/Y __dut__.__uuf__._1573_/A
+ __dut__.__uuf__._1988_/B VGND VGND VPWR VPWR __dut__.__uuf__._1984_/X sky130_fd_sc_hd__o22a_4
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0982_ __dut__._0982_/A __dut__._1907_/Q VGND VGND VPWR VPWR __dut__._0982_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1418_ __dut__.__uuf__._1418_/A VGND VGND VPWR VPWR __dut__.__uuf__._1418_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_78_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1697__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1603_ __dut__._1767_/A1 __dut__._1601_/X __dut__._1602_/X VGND VGND VPWR
+ VPWR __dut__._1804_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1349_ __dut__.__uuf__._1400_/A VGND VGND VPWR VPWR __dut__.__uuf__._1349_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1534_ rst VGND VGND VPWR VPWR __dut__._1534_/Y sky130_fd_sc_hd__inv_2
X__dut__._1465_ rst VGND VGND VPWR VPWR __dut__._1465_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1396_ __dut__._1408_/A prod[63] VGND VGND VPWR VPWR __dut__._1396_/X sky130_fd_sc_hd__and2_4
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1442__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1074__A __dut__.__uuf__._1551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1621__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_275_ _314_/CLK _275_/D VGND VGND VPWR VPWR _275_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1352__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_0_0___dut__.__uuf__.__clk_source__ clkbuf_4_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2065_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_87_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1203_ __dut__.__uuf__._1198_/X __dut__.__uuf__._1195_/X prod[21]
+ prod[22] __dut__.__uuf__._1191_/X VGND VGND VPWR VPWR __dut__._1311_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._2183_ __dut__.__uuf__._2194_/CLK __dut__._1355_/X __dut__.__uuf__._1137_/X
+ VGND VGND VPWR VPWR prod[43] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1527__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1134_ __dut__.__uuf__._1144_/A VGND VGND VPWR VPWR __dut__.__uuf__._1134_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1065_ __dut__.__uuf__._1328_/A VGND VGND VPWR VPWR __dut__.__uuf__._1314_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_67_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1250_ __dut__._1408_/A __dut__._1250_/B VGND VGND VPWR VPWR __dut__._1250_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1262__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1181_ __dut__._1193_/A1 __dut__._1181_/A2 __dut__._1180_/X VGND VGND VPWR
+ VPWR __dut__._1181_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2144__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1603__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1967_ __dut__.__uuf__._1961_/Y __dut__.__uuf__._1962_/Y __dut__.__uuf__._1961_/Y
+ __dut__.__uuf__._1962_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1968_/C sky130_fd_sc_hd__a2bb2o_4
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1898_ __dut__._0873_/X VGND VGND VPWR VPWR __dut__.__uuf__._1903_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_11_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpsn_inst_psn_buff_92 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1349_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_70 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1049_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_3_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_81 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1767_/A1
+ sky130_fd_sc_hd__buf_8
X__dut__._0965_ __dut__._0967_/A1 prod[14] __dut__._0964_/X VGND VGND VPWR VPWR __dut__._1899_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0896_ __dut__._1378_/A __dut__._1864_/Q VGND VGND VPWR VPWR __dut__._0896_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1437__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1517_ rst VGND VGND VPWR VPWR __dut__._1517_/Y sky130_fd_sc_hd__inv_2
X__dut__._1448_ rst VGND VGND VPWR VPWR __dut__._1448_/Y sky130_fd_sc_hd__inv_2
X__dut__._1379_ __dut__._1383_/A1 __dut__._1379_/A2 __dut__._1378_/X VGND VGND VPWR
+ VPWR __dut__._1379_/X sky130_fd_sc_hd__a21o_4
XFILLER_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_258_ _306_/CLK _258_/D VGND VGND VPWR VPWR _258_/Q sky130_fd_sc_hd__dfxtp_4
X_189_ _264_/Q _191_/B VGND VGND VPWR VPWR _263_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2017__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_161_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1821_ __dut__.__uuf__._1818_/Y __dut__.__uuf__._1819_/Y __dut__.__uuf__._1798_/X
+ __dut__.__uuf__._1825_/B VGND VGND VPWR VPWR __dut__.__uuf__._1821_/X sky130_fd_sc_hd__o22a_4
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1752_ __dut__._1042_/B VGND VGND VPWR VPWR __dut__.__uuf__._1752_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1683_ __dut__._1018_/B VGND VGND VPWR VPWR __dut__.__uuf__._1683_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_20_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2166_ __dut__.__uuf__._2169_/CLK __dut__._1321_/X __dut__.__uuf__._1187_/X
+ VGND VGND VPWR VPWR prod[26] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1117_ __dut__.__uuf__._1175_/A VGND VGND VPWR VPWR __dut__.__uuf__._1117_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0875__A2 __dut__._0873_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2097_ __dut__.__uuf__._2097_/CLK __dut__._1183_/X __dut__.__uuf__._1479_/X
+ VGND VGND VPWR VPWR __dut__._1184_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._1302_ __dut__._1302_/A prod[16] VGND VGND VPWR VPWR __dut__._1302_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1048_ __dut__.__uuf__._2008_/A VGND VGND VPWR VPWR __dut__.__uuf__._1063_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1233_ __dut__._1787_/A1 __dut__._1233_/A2 __dut__._1232_/X VGND VGND VPWR
+ VPWR __dut__._1233_/X sky130_fd_sc_hd__a21o_4
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1720__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1164_ __dut__._1766_/A __dut__._1164_/B VGND VGND VPWR VPWR __dut__._1164_/X
+ sky130_fd_sc_hd__and2_4
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1095_ __dut__._1129_/A1 __dut__._1095_/A2 __dut__._1094_/X VGND VGND VPWR
+ VPWR __dut__._1095_/X sky130_fd_sc_hd__a21o_4
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._0948_ __dut__._1770_/A __dut__._1890_/Q VGND VGND VPWR VPWR __dut__._0948_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0879_ __dut__._1409_/A1 prod[36] __dut__._0878_/X VGND VGND VPWR VPWR __dut__._1856_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_3_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2020_ __dut__.__uuf__._2049_/CLK __dut__._1029_/X __dut__.__uuf__._1642_/X
+ VGND VGND VPWR VPWR __dut__._1030_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_57_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__270__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1540__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1804_ __dut__.__uuf__._1804_/A __dut__.__uuf__._1804_/B __dut__.__uuf__._1804_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1806_/B sky130_fd_sc_hd__or3_4
XFILLER_21_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1735_ __dut__.__uuf__._1731_/Y __dut__.__uuf__._1732_/Y __dut__.__uuf__._1721_/X
+ __dut__.__uuf__._1734_/X VGND VGND VPWR VPWR __dut__.__uuf__._1736_/A sky130_fd_sc_hd__a211o_4
X__dut__.__uuf__._1666_ __dut__.__uuf__._1781_/A VGND VGND VPWR VPWR __dut__.__uuf__._1717_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1597_ __dut__.__uuf__._1599_/A VGND VGND VPWR VPWR __dut__.__uuf__._1597_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1851_ __dut__._1410_/B __dut__._1851_/D __dut__._1478_/Y VGND VGND VPWR
+ VPWR __dut__._1851_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1782_ __dut__._1786_/A __dut__._1848_/Q VGND VGND VPWR VPWR __dut__._1782_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2149_ __dut__.__uuf__._2169_/CLK __dut__._1287_/X __dut__.__uuf__._1237_/X
+ VGND VGND VPWR VPWR prod[9] sky130_fd_sc_hd__dfrtp_4
XFILLER_75_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_62_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1216_ __dut__._1786_/A __dut__._1216_/B VGND VGND VPWR VPWR __dut__._1216_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1450__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1147_ __dut__._1647_/A1 __dut__._1147_/A2 __dut__._1146_/X VGND VGND VPWR
+ VPWR __dut__._1147_/X sky130_fd_sc_hd__a21o_4
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1078_ __dut__._1078_/A __dut__._1078_/B VGND VGND VPWR VPWR __dut__._1078_/X
+ sky130_fd_sc_hd__and2_4
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2205__CLK __dut__.__uuf__._2210_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_124_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1360__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_10_0_tck clkbuf_3_5_0_tck/X VGND VGND VPWR VPWR __dut__._1883_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1520_ __dut__._1697_/X __dut__.__uuf__._1515_/X __dut__._1168_/B
+ __dut__.__uuf__._1516_/X VGND VGND VPWR VPWR __dut__.__uuf__._1520_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__._1817__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1720__A __dut__.__uuf__._1720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1451_ __dut__.__uuf__._1566_/A VGND VGND VPWR VPWR __dut__.__uuf__._1451_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1382_ __dut__.__uuf__._1381_/Y __dut__.__uuf__._1375_/X __dut__.__uuf__._1376_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1382_/X sky130_fd_sc_hd__o21a_4
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1535__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2003_ __dut__.__uuf__._2003_/A __dut__.__uuf__._2003_/B __dut__.__uuf__._2003_/C
+ VGND VGND VPWR VPWR __dut__._1131_/A2 sky130_fd_sc_hd__and3_4
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1001_ __dut__._1339_/A1 prod[32] __dut__._1000_/X VGND VGND VPWR VPWR __dut__._1917_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA__303__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1718_ __dut__._1030_/B VGND VGND VPWR VPWR __dut__.__uuf__._1718_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1649_ __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR __dut__.__uuf__._1654_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1903_ clkbuf_4_9_0_tck/X __dut__._1903_/D __dut__._1426_/Y VGND VGND VPWR
+ VPWR __dut__._1903_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1834_ __dut__._1410_/B __dut__._1834_/D __dut__._1495_/Y VGND VGND VPWR
+ VPWR __dut__._1834_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1765_ __dut__._1543_/Y mc[5] __dut__._1764_/X VGND VGND VPWR VPWR __dut__._1765_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1696_ __dut__._1788_/A __dut__._1828_/Q VGND VGND VPWR VPWR __dut__._1696_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1445__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1077__A __dut__.__uuf__._1450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__.__uuf__._1081__A3 prod[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1503_ __dut__.__uuf__._1487_/X __dut__.__uuf__._1483_/X __dut__._1174_/B
+ __dut__.__uuf__._1493_/X __dut__.__uuf__._1502_/X VGND VGND VPWR VPWR __dut__._1173_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__.__uuf__._1450__A __dut__.__uuf__._1450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1434_ __dut__.__uuf__._1433_/Y __dut__.__uuf__._1425_/X __dut__.__uuf__._1324_/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._1434_/X sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._1173__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1365_ __dut__.__uuf__._1380_/A VGND VGND VPWR VPWR __dut__.__uuf__._1365_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_89_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1550_ __dut__._1766_/A __dut__._1854_/Q VGND VGND VPWR VPWR __dut__._1550_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1296_ __dut__.__uuf__._1720_/A VGND VGND VPWR VPWR __dut__.__uuf__._1400_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_85_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1481_ rst VGND VGND VPWR VPWR __dut__._1481_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_291_ _313_/CLK _291_/D trst VGND VGND VPWR VPWR _291_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_25_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1817_ clkbuf_4_5_0_tck/X __dut__._1817_/D __dut__._1512_/Y VGND VGND VPWR
+ VPWR __dut__._1817_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._0911__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1748_ __dut__._1788_/A __dut__._1841_/Q VGND VGND VPWR VPWR __dut__._1748_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1679_ __dut__._1679_/A1 __dut__._1677_/X __dut__._1678_/X VGND VGND VPWR
+ VPWR __dut__._1823_/D sky130_fd_sc_hd__a21o_4
XANTENNA__296__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1150_ __dut__.__uuf__._1138_/X __dut__.__uuf__._1149_/X prod[39]
+ prod[40] __dut__.__uuf__._1145_/X VGND VGND VPWR VPWR __dut__._1347_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_101_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1081_ __dut__.__uuf__._1075_/X __dut__.__uuf__._2003_/A prod[62]
+ prod[63] __dut__.__uuf__._1069_/X VGND VGND VPWR VPWR __dut__._1393_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1983_ __dut__._1589_/X VGND VGND VPWR VPWR __dut__.__uuf__._1988_/B
+ sky130_fd_sc_hd__inv_2
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._0981_ __dut__._0981_/A1 prod[22] __dut__._0980_/X VGND VGND VPWR VPWR __dut__._1907_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2073__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1417_ __dut__.__uuf__._1405_/X __dut__.__uuf__._1415_/X __dut__._1212_/B
+ __dut__.__uuf__._1416_/X VGND VGND VPWR VPWR __dut__._1211_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1602_ __dut__._1766_/A __dut__._1803_/Q VGND VGND VPWR VPWR __dut__._1602_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1697__A2 mp[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1348_ __dut__._1240_/B VGND VGND VPWR VPWR __dut__.__uuf__._1348_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1533_ rst VGND VGND VPWR VPWR __dut__._1533_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1279_ __dut__.__uuf__._1288_/A VGND VGND VPWR VPWR __dut__.__uuf__._1279_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1464_ rst VGND VGND VPWR VPWR __dut__._1464_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1395_ __dut__._1395_/A1 __dut__._1395_/A2 __dut__._1394_/X VGND VGND VPWR
+ VPWR __dut__._1395_/X sky130_fd_sc_hd__a21o_4
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1621__A2 mc[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_274_ _314_/CLK _274_/D VGND VGND VPWR VPWR _274_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1202_ __dut__.__uuf__._1204_/A VGND VGND VPWR VPWR __dut__.__uuf__._1202_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2182_ __dut__.__uuf__._2194_/CLK __dut__._1353_/X __dut__.__uuf__._1140_/X
+ VGND VGND VPWR VPWR prod[42] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1133_ __dut__.__uuf__._1162_/A VGND VGND VPWR VPWR __dut__.__uuf__._1144_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1064_ __dut__._1400_/B __dut__._1398_/B VGND VGND VPWR VPWR __dut__.__uuf__._1064_/X
+ sky130_fd_sc_hd__or2_4
XANTENNA___dut__._1543__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1180_ __dut__._1180_/A __dut__._1180_/B VGND VGND VPWR VPWR __dut__._1180_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1966_ __dut__.__uuf__._1966_/A VGND VGND VPWR VPWR __dut__._1117_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1897_ __dut__._1088_/B VGND VGND VPWR VPWR __dut__.__uuf__._1897_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_7_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1367__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_71 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1057_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1119__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_60 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1165_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1718__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_82 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1719_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._0964_ __dut__._1324_/A __dut__._1898_/Q VGND VGND VPWR VPWR __dut__._0964_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_93 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1395_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._0895_ __dut__._1383_/A1 prod[44] __dut__._0894_/X VGND VGND VPWR VPWR __dut__._1864_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_92_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_10_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2206_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__._1516_ rst VGND VGND VPWR VPWR __dut__._1516_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1453__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1085__A __dut__.__uuf__._1100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1447_ rst VGND VGND VPWR VPWR __dut__._1447_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1378_ __dut__._1378_/A prod[54] VGND VGND VPWR VPWR __dut__._1378_/X sky130_fd_sc_hd__and2_4
XFILLER_34_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_257_ _306_/CLK _257_/D VGND VGND VPWR VPWR _258_/D sky130_fd_sc_hd__dfxtp_4
X_188_ _265_/Q _191_/B VGND VGND VPWR VPWR _264_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1628__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1850__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_154_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1820_ __dut__._1573_/X VGND VGND VPWR VPWR __dut__.__uuf__._1825_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1597__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1751_ __dut__.__uuf__._1773_/A __dut__.__uuf__._1751_/B __dut__.__uuf__._1751_/C
+ VGND VGND VPWR VPWR __dut__._1035_/A2 sky130_fd_sc_hd__and3_4
X__dut__.__uuf__._1682_ __dut__.__uuf__._1717_/A __dut__.__uuf__._1682_/B __dut__.__uuf__._1682_/C
+ VGND VGND VPWR VPWR __dut__._1011_/A2 sky130_fd_sc_hd__and3_4
XANTENNA___dut__._1538__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2165_ __dut__.__uuf__._2169_/CLK __dut__._1319_/X __dut__.__uuf__._1189_/X
+ VGND VGND VPWR VPWR prod[25] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._2111__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1116_ __dut__.__uuf__._1190_/A VGND VGND VPWR VPWR __dut__.__uuf__._1175_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2096_ __dut__.__uuf__._2097_/CLK __dut__._1181_/X __dut__.__uuf__._1482_/X
+ VGND VGND VPWR VPWR __dut__._1182_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._1301_ __dut__._1301_/A1 __dut__._1301_/A2 __dut__._1300_/X VGND VGND VPWR
+ VPWR __dut__._1301_/X sky130_fd_sc_hd__a21o_4
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1047_ __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR __dut__.__uuf__._2008_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_71_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1232_ __dut__._1786_/A __dut__._1232_/B VGND VGND VPWR VPWR __dut__._1232_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1163_ __dut__._1163_/A1 __dut__._1163_/A2 __dut__._1162_/X VGND VGND VPWR
+ VPWR __dut__._1163_/X sky130_fd_sc_hd__a21o_4
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1949_ __dut__.__uuf__._1936_/X __dut__.__uuf__._1948_/B __dut__.__uuf__._1948_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1950_/C sky130_fd_sc_hd__o21ai_4
X__dut__._1094_ __dut__._1094_/A __dut__._1094_/B VGND VGND VPWR VPWR __dut__._1094_/X
+ sky130_fd_sc_hd__and2_4
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1873__CLK __dut__._1917_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1448__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0947_ __dut__._0947_/A1 prod[5] __dut__._0946_/X VGND VGND VPWR VPWR __dut__._1890_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0878_ __dut__._1408_/A __dut__._1855_/Q VGND VGND VPWR VPWR __dut__._0878_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1579__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_309_ _314_/CLK _309_/D trst VGND VGND VPWR VPWR _309_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1358__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1896__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1803_ __dut__.__uuf__._1796_/Y __dut__.__uuf__._1797_/Y __dut__.__uuf__._1796_/Y
+ __dut__.__uuf__._1797_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1804_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1734_ __dut__.__uuf__._1731_/Y __dut__.__uuf__._1732_/Y __dut__.__uuf__._1686_/X
+ __dut__.__uuf__._1738_/B VGND VGND VPWR VPWR __dut__.__uuf__._1734_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1665_ __dut__.__uuf__._1665_/A VGND VGND VPWR VPWR __dut__._1009_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1596_ __dut__.__uuf__._1599_/A VGND VGND VPWR VPWR __dut__.__uuf__._1596_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1850_ _194_/A __dut__._1850_/D __dut__._1479_/Y VGND VGND VPWR VPWR __dut__._1850_/Q
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1268__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1781_ __dut__._1543_/Y mp[31] __dut__._1780_/X VGND VGND VPWR VPWR __dut__._1781_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._0900__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2148_ __dut__.__uuf__._2169_/CLK __dut__._1285_/X __dut__.__uuf__._1241_/X
+ VGND VGND VPWR VPWR prod[8] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2079_ __dut__.__uuf__._2107_/CLK __dut__._1147_/X __dut__.__uuf__._1555_/X
+ VGND VGND VPWR VPWR __dut__._1148_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_55_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1215_ __dut__._1787_/A1 __dut__._1215_/A2 __dut__._1214_/X VGND VGND VPWR
+ VPWR __dut__._1215_/X sky130_fd_sc_hd__a21o_4
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1146_ __dut__._1146_/A __dut__._1146_/B VGND VGND VPWR VPWR __dut__._1146_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0___dut__.__uuf__.__clk_source__ clkbuf_4_9_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2208_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__._1077_ __dut__._1129_/A1 __dut__._1077_/A2 __dut__._1076_/X VGND VGND VPWR
+ VPWR __dut__._1077_/X sky130_fd_sc_hd__a21o_4
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1733__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0___dut__.__uuf__.__clk_source__ clkbuf_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR clkbuf_2_3_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__157__A tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_117_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1450_ __dut__.__uuf__._1450_/A VGND VGND VPWR VPWR __dut__.__uuf__._1566_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1381_ __dut__._1228_/B VGND VGND VPWR VPWR __dut__.__uuf__._1381_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_89_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2002_ __dut__.__uuf__._1692_/A __dut__.__uuf__._2001_/B __dut__.__uuf__._2001_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2003_/C sky130_fd_sc_hd__o21ai_4
XFILLER_85_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1000_ __dut__._1378_/A __dut__._1916_/Q VGND VGND VPWR VPWR __dut__._1000_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1270__B prod[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1717_ __dut__.__uuf__._1717_/A __dut__.__uuf__._1717_/B __dut__.__uuf__._1717_/C
+ VGND VGND VPWR VPWR __dut__._1023_/A2 sky130_fd_sc_hd__and3_4
XFILLER_5_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1648_ __dut__.__uuf__._1648_/A VGND VGND VPWR VPWR __dut__.__uuf__._1648_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1902_ __dut__._1902_/CLK __dut__._1902_/D __dut__._1427_/Y VGND VGND VPWR
+ VPWR __dut__._1902_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1833_ clkbuf_4_7_0_tck/X __dut__._1833_/D __dut__._1496_/Y VGND VGND VPWR
+ VPWR __dut__._1833_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1911__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1579_ __dut__.__uuf__._1580_/A VGND VGND VPWR VPWR __dut__.__uuf__._1579_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1764_ __dut__._1788_/A __dut__._1845_/Q VGND VGND VPWR VPWR __dut__._1764_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1695_ __dut__._1719_/A1 __dut__._1693_/X __dut__._1694_/X VGND VGND VPWR
+ VPWR __dut__._1827_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1726__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1461__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1129_ __dut__._1129_/A1 __dut__._1129_/A2 __dut__._1128_/X VGND VGND VPWR
+ VPWR __dut__._1129_/X sky130_fd_sc_hd__a21o_4
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__260__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1636__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1502_ __dut__._1713_/X __dut__.__uuf__._1494_/X __dut__._1176_/B
+ __dut__.__uuf__._1495_/X VGND VGND VPWR VPWR __dut__.__uuf__._1502_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1433_ __dut__._1206_/B VGND VGND VPWR VPWR __dut__.__uuf__._1433_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1364_ __dut__.__uuf__._1363_/Y __dut__.__uuf__._1349_/X __dut__.__uuf__._1350_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1364_/X sky130_fd_sc_hd__o21a_4
XFILLER_89_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1546__A tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1295_ __dut__.__uuf__._1295_/A VGND VGND VPWR VPWR __dut__.__uuf__._1720_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1480_ rst VGND VGND VPWR VPWR __dut__._1480_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_290_ _290_/CLK _290_/D VGND VGND VPWR VPWR _290_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__283__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_18_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1816_ clkbuf_4_6_0_tck/X __dut__._1816_/D __dut__._1513_/Y VGND VGND VPWR
+ VPWR __dut__._1816_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1456__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1747_ __dut__._1759_/A1 __dut__._1745_/X __dut__._1746_/X VGND VGND VPWR
+ VPWR __dut__._1840_/D sky130_fd_sc_hd__a21o_4
X__dut__._1678_ __dut__._1678_/A __dut__._1812_/Q VGND VGND VPWR VPWR __dut__._1678_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1807__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__.__uuf__._1551__A __dut__.__uuf__._1551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1366__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1080_ __dut__.__uuf__._1084_/A VGND VGND VPWR VPWR __dut__.__uuf__._1080_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1982_ __dut__._1120_/B VGND VGND VPWR VPWR __dut__.__uuf__._1982_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1091__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0980_ __dut__._1404_/A __dut__._1906_/Q VGND VGND VPWR VPWR __dut__._0980_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1416_ __dut__.__uuf__._1416_/A VGND VGND VPWR VPWR __dut__.__uuf__._1416_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1601_ __dut__._1543_/Y mc[22] __dut__._1600_/X VGND VGND VPWR VPWR __dut__._1601_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1347_ __dut__.__uuf__._1367_/A VGND VGND VPWR VPWR __dut__.__uuf__._1347_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1532_ rst VGND VGND VPWR VPWR __dut__._1532_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1278_ __dut__.__uuf__._1274_/X __dut__.__uuf__._1277_/X __dut__._1266_/B
+ __dut__.__uuf__._1274_/X VGND VGND VPWR VPWR __dut__._1265_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1463_ rst VGND VGND VPWR VPWR __dut__._1463_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1394_ __dut__._1542_/A prod[62] VGND VGND VPWR VPWR __dut__._1394_/X sky130_fd_sc_hd__and2_4
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_273_ _314_/CLK _273_/D VGND VGND VPWR VPWR _273_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__.__uuf__._1371__A __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1186__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1073__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1201_ __dut__.__uuf__._1198_/X __dut__.__uuf__._1195_/X prod[22]
+ prod[23] __dut__.__uuf__._1191_/X VGND VGND VPWR VPWR __dut__._1313_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1096__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2181_ __dut__.__uuf__._2200_/CLK __dut__._1351_/X __dut__.__uuf__._1142_/X
+ VGND VGND VPWR VPWR prod[41] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1132_ __dut__.__uuf__._1124_/X __dut__.__uuf__._1121_/X prod[45]
+ prod[46] __dut__.__uuf__._1131_/X VGND VGND VPWR VPWR __dut__._1359_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1063_ __dut__.__uuf__._1063_/A VGND VGND VPWR VPWR __dut__.__uuf__._1063_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1965_ __dut__.__uuf__._1961_/Y __dut__.__uuf__._1962_/Y __dut__.__uuf__._1941_/X
+ __dut__.__uuf__._1964_/X VGND VGND VPWR VPWR __dut__.__uuf__._1966_/A sky130_fd_sc_hd__a211o_4
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1896_ __dut__._1094_/B VGND VGND VPWR VPWR __dut__.__uuf__._1896_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0963_ __dut__._0967_/A1 prod[13] __dut__._0962_/X VGND VGND VPWR VPWR __dut__._1898_/D
+ sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_72 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1055_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_61 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1163_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_50 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0949_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_83 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1289_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._0894_ __dut__._1378_/A __dut__._1863_/Q VGND VGND VPWR VPWR __dut__._0894_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_94 _244_/X VGND VGND VPWR VPWR __dut__._1678_/A sky130_fd_sc_hd__buf_8
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0___dut__.__uuf__.__clk_source__ clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_5_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
X__dut__._1515_ rst VGND VGND VPWR VPWR __dut__._1515_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1734__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1446_ rst VGND VGND VPWR VPWR __dut__._1446_/Y sky130_fd_sc_hd__inv_2
X__dut__._1377_ __dut__._1383_/A1 __dut__._1377_/A2 __dut__._1376_/X VGND VGND VPWR
+ VPWR __dut__._1377_/X sky130_fd_sc_hd__a21o_4
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_256_ _306_/CLK _256_/D VGND VGND VPWR VPWR _257_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_6_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_187_ _266_/Q _187_/B VGND VGND VPWR VPWR _265_/D sky130_fd_sc_hd__or2_4
XFILLER_96_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0869__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1644__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_147_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1750_ __dut__.__uuf__._1715_/X __dut__.__uuf__._1749_/B __dut__.__uuf__._1749_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1751_/C sky130_fd_sc_hd__o21ai_4
XANTENNA___dut__._1597__A2 mc[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1681_ __dut__.__uuf__._1573_/X __dut__.__uuf__._1680_/B __dut__.__uuf__._1680_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1682_/C sky130_fd_sc_hd__o21ai_4
X__dut__.__uuf__._2164_ __dut__.__uuf__._2164_/CLK __dut__._1317_/X __dut__.__uuf__._1194_/X
+ VGND VGND VPWR VPWR prod[24] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1115_ __dut__.__uuf__._1115_/A VGND VGND VPWR VPWR __dut__.__uuf__._1115_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1554__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1300_ __dut__._1324_/A prod[15] VGND VGND VPWR VPWR __dut__._1300_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._2095_ __dut__.__uuf__._2107_/CLK __dut__._1179_/X __dut__.__uuf__._1486_/X
+ VGND VGND VPWR VPWR __dut__._1180_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1046_ __dut__.__uuf__._1102_/A VGND VGND VPWR VPWR __dut__.__uuf__._1612_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1231_ __dut__._1787_/A1 __dut__._1231_/A2 __dut__._1230_/X VGND VGND VPWR
+ VPWR __dut__._1231_/X sky130_fd_sc_hd__a21o_4
X__dut__._1162_ __dut__._1766_/A __dut__._1162_/B VGND VGND VPWR VPWR __dut__._1162_/X
+ sky130_fd_sc_hd__and2_4
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1948_ __dut__.__uuf__._1968_/A __dut__.__uuf__._1948_/B __dut__.__uuf__._1948_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1950_/B sky130_fd_sc_hd__or3_4
X__dut__._1093_ __dut__._1129_/A1 __dut__._1093_/A2 __dut__._1092_/X VGND VGND VPWR
+ VPWR __dut__._1093_/X sky130_fd_sc_hd__a21o_4
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1879_ __dut__.__uuf__._1873_/Y __dut__.__uuf__._1874_/Y __dut__.__uuf__._1873_/Y
+ __dut__.__uuf__._1874_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1880_/C sky130_fd_sc_hd__a2bb2o_4
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._0946_ __dut__._1770_/A __dut__._1889_/Q VGND VGND VPWR VPWR __dut__._0946_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_78_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._0877_ __dut__._0877_/A1 prod[35] __dut__._0876_/X VGND VGND VPWR VPWR __dut__._1855_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1464__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1429_ rst VGND VGND VPWR VPWR __dut__._1429_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_308_ _314_/CLK _308_/D trst VGND VGND VPWR VPWR _308_/Q sky130_fd_sc_hd__dfrtp_4
X_239_ _239_/A _302_/Q _239_/C VGND VGND VPWR VPWR _251_/D sky130_fd_sc_hd__or3_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1374__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1267__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1019__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1802_ __dut__.__uuf__._1802_/A VGND VGND VPWR VPWR __dut__._1057_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1733_ __dut__._1609_/X VGND VGND VPWR VPWR __dut__.__uuf__._1738_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1664_ __dut__.__uuf__._1658_/Y __dut__.__uuf__._1659_/Y __dut__.__uuf__._1660_/X
+ __dut__.__uuf__._1663_/X VGND VGND VPWR VPWR __dut__.__uuf__._1665_/A sky130_fd_sc_hd__a211o_4
X__dut__.__uuf__._1595_ __dut__.__uuf__._1599_/A VGND VGND VPWR VPWR __dut__.__uuf__._1595_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1780_ __dut__._1788_/A __dut__._1849_/Q VGND VGND VPWR VPWR __dut__._1780_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1909__A __dut__._0869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1284__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2147_ __dut__.__uuf__._2164_/CLK __dut__._1283_/X __dut__.__uuf__._1244_/X
+ VGND VGND VPWR VPWR prod[7] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2078_ __dut__.__uuf__._2107_/CLK __dut__._1145_/X __dut__.__uuf__._1559_/X
+ VGND VGND VPWR VPWR __dut__._1146_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1029_ __dut__.__uuf__._1029_/A __dut__.__uuf__._1029_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1061_/B sky130_fd_sc_hd__or2_4
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1840__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1214_ __dut__._1786_/A __dut__._1214_/B VGND VGND VPWR VPWR __dut__._1214_/X
+ sky130_fd_sc_hd__and2_4
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_48_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1145_ __dut__._1647_/A1 __dut__._1145_/A2 __dut__._1144_/X VGND VGND VPWR
+ VPWR __dut__._1145_/X sky130_fd_sc_hd__a21o_4
XFILLER_101_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1076_ __dut__._1678_/A __dut__._1076_/B VGND VGND VPWR VPWR __dut__._1076_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_12_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1459__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1733__A2 mp[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0929_ __dut__._1395_/A1 prod[61] __dut__._0928_/X VGND VGND VPWR VPWR __dut__._1881_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1249__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2101__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1380_ __dut__.__uuf__._1380_/A VGND VGND VPWR VPWR __dut__.__uuf__._1380_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2001_ __dut__.__uuf__._2001_/A __dut__.__uuf__._2001_/B __dut__.__uuf__._2001_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._2003_/B sky130_fd_sc_hd__or3_4
XANTENNA___dut__._1863__CLK __dut__._1917_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1716_ __dut__.__uuf__._1715_/X __dut__.__uuf__._1713_/B __dut__.__uuf__._1713_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1717_/C sky130_fd_sc_hd__o21ai_4
X__dut__.__uuf__._1647_ __dut__.__uuf__._1648_/A VGND VGND VPWR VPWR __dut__.__uuf__._1647_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1901_ __dut__._1902_/CLK __dut__._1901_/D __dut__._1428_/Y VGND VGND VPWR
+ VPWR __dut__._1901_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1832_ __dut__._1899_/CLK __dut__._1832_/D __dut__._1497_/Y VGND VGND VPWR
+ VPWR __dut__._1832_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1578_ __dut__.__uuf__._1580_/A VGND VGND VPWR VPWR __dut__.__uuf__._1578_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1763_ __dut__._1763_/A1 __dut__._1761_/X __dut__._1762_/X VGND VGND VPWR
+ VPWR __dut__._1844_/D sky130_fd_sc_hd__a21o_4
X__dut__._1694_ __dut__._1766_/A __dut__._1826_/Q VGND VGND VPWR VPWR __dut__._1694_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1742__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1128_ __dut__._1128_/A __dut__._1128_/B VGND VGND VPWR VPWR __dut__._1128_/X
+ sky130_fd_sc_hd__and2_4
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1059_ __dut__._1767_/A1 __dut__._1059_/A2 __dut__._1058_/X VGND VGND VPWR
+ VPWR __dut__._1059_/X sky130_fd_sc_hd__a21o_4
XFILLER_8_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1652__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1501_ __dut__.__uuf__._1508_/A VGND VGND VPWR VPWR __dut__.__uuf__._1501_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_2_2_0_tck_A clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1432_ __dut__.__uuf__._1442_/A VGND VGND VPWR VPWR __dut__.__uuf__._1432_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1363_ __dut__._1234_/B VGND VGND VPWR VPWR __dut__.__uuf__._1363_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1294_ __dut__._1260_/B VGND VGND VPWR VPWR __dut__.__uuf__._1294_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_58_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1562__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2147__CLK __dut__.__uuf__._2164_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1633__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0906__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1815_ clkbuf_4_6_0_tck/X __dut__._1815_/D __dut__._1514_/Y VGND VGND VPWR
+ VPWR __dut__._1815_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1746_ __dut__._1770_/A __dut__._1839_/Q VGND VGND VPWR VPWR __dut__._1746_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1677_ __dut__._1543_/Y mc[3] __dut__._1676_/X VGND VGND VPWR VPWR __dut__._1677_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_1_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1472__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1382__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1615__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1981_ __dut__._1126_/B VGND VGND VPWR VPWR __dut__.__uuf__._1981_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1901__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1415_ __dut__.__uuf__._1414_/Y __dut__.__uuf__._1400_/X __dut__.__uuf__._1401_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1415_/X sky130_fd_sc_hd__o21a_4
X__dut__._1600_ __dut__._1788_/A __dut__._1804_/Q VGND VGND VPWR VPWR __dut__._1600_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1276__B prod[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1346_ __dut__.__uuf__._1346_/A VGND VGND VPWR VPWR __dut__.__uuf__._1367_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1531_ rst VGND VGND VPWR VPWR __dut__._1531_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1277_ __dut__.__uuf__._1267_/Y __dut__.__uuf__._1276_/X __dut__.__uuf__._1271_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1277_/X sky130_fd_sc_hd__o21a_4
X__dut__._1462_ rst VGND VGND VPWR VPWR __dut__._1462_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1393_ __dut__._1395_/A1 __dut__._1393_/A2 __dut__._1392_/X VGND VGND VPWR
+ VPWR __dut__._1393_/X sky130_fd_sc_hd__a21o_4
XFILLER_85_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_0 __dut__._1542_/Y VGND VGND VPWR VPWR psn_inst_psn_buff_9/A sky130_fd_sc_hd__buf_8
X_272_ _314_/CLK _272_/D VGND VGND VPWR VPWR _272_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_psn_inst_psn_buff_30_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1467__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1729_ __dut__._1543_/Y mp[19] __dut__._1728_/X VGND VGND VPWR VPWR __dut__._1729_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2180_ __dut__.__uuf__._2200_/CLK __dut__._1349_/X __dut__.__uuf__._1144_/X
+ VGND VGND VPWR VPWR prod[40] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1200_ __dut__.__uuf__._1204_/A VGND VGND VPWR VPWR __dut__.__uuf__._1200_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._1131_ __dut__.__uuf__._1175_/A VGND VGND VPWR VPWR __dut__.__uuf__._1131_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1062_ __dut__.__uuf__._1031_/A __dut__.__uuf__._1061_/Y __dut__.__uuf__._1054_/X
+ __dut__._1402_/B __dut__.__uuf__._1043_/X VGND VGND VPWR VPWR __dut__._1401_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA__273__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1964_ __dut__.__uuf__._1961_/Y __dut__.__uuf__._1962_/Y __dut__.__uuf__._1573_/A
+ __dut__.__uuf__._1968_/B VGND VGND VPWR VPWR __dut__.__uuf__._1964_/X sky130_fd_sc_hd__o22a_4
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1472__A __dut__.__uuf__._1536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1895_ __dut__.__uuf__._1938_/A __dut__.__uuf__._1895_/B __dut__.__uuf__._1895_/C
+ VGND VGND VPWR VPWR __dut__._1087_/A2 sky130_fd_sc_hd__and3_4
X__dut__._0962_ __dut__._1324_/A __dut__._1897_/Q VGND VGND VPWR VPWR __dut__._0962_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_40 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._0967_/A1
+ sky130_fd_sc_hd__buf_4
Xpsn_inst_psn_buff_73 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1053_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_62 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1161_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_51 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1187_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._0893_ __dut__._1383_/A1 prod[43] __dut__._0892_/X VGND VGND VPWR VPWR __dut__._1863_/D
+ sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_95 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1008_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_84 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR psn_inst_psn_buff_88/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1329_ __dut__.__uuf__._1380_/A VGND VGND VPWR VPWR __dut__.__uuf__._1329_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1514_ rst VGND VGND VPWR VPWR __dut__._1514_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_78_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1445_ rst VGND VGND VPWR VPWR __dut__._1445_/Y sky130_fd_sc_hd__inv_2
X__dut__._1376_ __dut__._1378_/A prod[53] VGND VGND VPWR VPWR __dut__._1376_/X sky130_fd_sc_hd__and2_4
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1750__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_255_ _306_/CLK tms VGND VGND VPWR VPWR _256_/D sky130_fd_sc_hd__dfxtp_4
X_186_ _267_/Q _187_/B VGND VGND VPWR VPWR _266_/D sky130_fd_sc_hd__or2_4
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0869__A2 mc[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2208__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1660__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1680_ __dut__.__uuf__._1692_/A __dut__.__uuf__._1680_/B __dut__.__uuf__._1680_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1682_/B sky130_fd_sc_hd__or3_4
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._2163_ __dut__.__uuf__._2164_/CLK __dut__._1315_/X __dut__.__uuf__._1197_/X
+ VGND VGND VPWR VPWR prod[23] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1114_ __dut__.__uuf__._1109_/X __dut__.__uuf__._1106_/X prod[51]
+ prod[52] __dut__.__uuf__._1100_/X VGND VGND VPWR VPWR __dut__._1371_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_87_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2094_ __dut__.__uuf__._2107_/CLK __dut__._1177_/X __dut__.__uuf__._1492_/X
+ VGND VGND VPWR VPWR __dut__._1178_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1045_ rst VGND VGND VPWR VPWR __dut__.__uuf__._1102_/A sky130_fd_sc_hd__inv_2
X__dut__._1230_ __dut__._1786_/A __dut__._1230_/B VGND VGND VPWR VPWR __dut__._1230_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1570__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1161_ __dut__._1161_/A1 __dut__._1161_/A2 __dut__._1160_/X VGND VGND VPWR
+ VPWR __dut__._1161_/X sky130_fd_sc_hd__a21o_4
XFILLER_36_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1947_ __dut__.__uuf__._1939_/Y __dut__.__uuf__._1940_/Y __dut__.__uuf__._1939_/Y
+ __dut__.__uuf__._1940_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1948_/C sky130_fd_sc_hd__a2bb2o_4
X__dut__._1092_ __dut__._1094_/A __dut__._1092_/B VGND VGND VPWR VPWR __dut__._1092_/X
+ sky130_fd_sc_hd__and2_4
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1878_ __dut__.__uuf__._1878_/A VGND VGND VPWR VPWR __dut__._1085_/A2
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._0914__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1930__A __dut__._1789_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0945_ __dut__._0945_/A1 prod[4] __dut__._0944_/X VGND VGND VPWR VPWR __dut__._1889_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0876_ __dut__._0876_/A __dut__._1919_/Q VGND VGND VPWR VPWR __dut__._0876_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1428_ rst VGND VGND VPWR VPWR __dut__._1428_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1480__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1359_ __dut__._1383_/A1 __dut__._1359_/A2 __dut__._1358_/X VGND VGND VPWR
+ VPWR __dut__._1359_/X sky130_fd_sc_hd__a21o_4
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_307_ _194_/A _307_/D trst VGND VGND VPWR VPWR _307_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_238_ _238_/A _238_/B _300_/Q _238_/D VGND VGND VPWR VPWR _239_/C sky130_fd_sc_hd__and4_4
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_169_ _281_/Q _173_/B VGND VGND VPWR VPWR _280_/D sky130_fd_sc_hd__and2_4
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2030__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_84_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1390__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__311__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1801_ __dut__.__uuf__._1796_/Y __dut__.__uuf__._1797_/Y __dut__.__uuf__._1776_/X
+ __dut__.__uuf__._1800_/X VGND VGND VPWR VPWR __dut__.__uuf__._1802_/A sky130_fd_sc_hd__a211o_4
X__dut__.__uuf__._1732_ __dut__._1028_/B VGND VGND VPWR VPWR __dut__.__uuf__._1732_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1663_ __dut__.__uuf__._1658_/Y __dut__.__uuf__._1659_/Y __dut__.__uuf__._2001_/A
+ __dut__.__uuf__._1670_/B VGND VGND VPWR VPWR __dut__.__uuf__._1663_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__._1792__CLK __dut__._1410_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1594_ __dut__.__uuf__._1606_/A VGND VGND VPWR VPWR __dut__.__uuf__._1599_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2146_ __dut__.__uuf__._2164_/CLK __dut__._1281_/X __dut__.__uuf__._1246_/X
+ VGND VGND VPWR VPWR prod[6] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2077_ __dut__.__uuf__._2107_/CLK __dut__._1143_/X __dut__.__uuf__._1562_/X
+ VGND VGND VPWR VPWR __dut__._1144_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1028_ __dut__._1398_/B VGND VGND VPWR VPWR __dut__.__uuf__._1029_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1213_ __dut__._1787_/A1 __dut__._1213_/A2 __dut__._1212_/X VGND VGND VPWR
+ VPWR __dut__._1213_/X sky130_fd_sc_hd__a21o_4
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1144_ __dut__._1144_/A __dut__._1144_/B VGND VGND VPWR VPWR __dut__._1144_/X
+ sky130_fd_sc_hd__and2_4
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1075_ __dut__._1075_/A1 __dut__._1075_/A2 __dut__._1074_/X VGND VGND VPWR
+ VPWR __dut__._1075_/X sky130_fd_sc_hd__a21o_4
XFILLER_24_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._0928_ __dut__._1542_/A __dut__._1880_/Q VGND VGND VPWR VPWR __dut__._0928_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1475__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2000_ __dut__.__uuf__._1994_/Y __dut__.__uuf__._1995_/Y __dut__.__uuf__._1994_/Y
+ __dut__.__uuf__._1995_/Y VGND VGND VPWR VPWR __dut__.__uuf__._2001_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1715_ __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR __dut__.__uuf__._1715_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1646_ __dut__.__uuf__._1648_/A VGND VGND VPWR VPWR __dut__.__uuf__._1646_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2076__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1900_ __dut__._1902_/CLK __dut__._1900_/D __dut__._1429_/Y VGND VGND VPWR
+ VPWR __dut__._1900_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1831_ __dut__._1899_/CLK __dut__._1831_/D __dut__._1498_/Y VGND VGND VPWR
+ VPWR __dut__._1831_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1577_ __dut__.__uuf__._1580_/A VGND VGND VPWR VPWR __dut__.__uuf__._1577_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._0923__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1762_ __dut__._1770_/A __dut__._1843_/Q VGND VGND VPWR VPWR __dut__._1762_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1693_ __dut__._1543_/Y mp[11] __dut__._1692_/X VGND VGND VPWR VPWR __dut__._1693_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2129_ __dut__.__uuf__._2206_/CLK __dut__._1247_/X __dut__.__uuf__._1321_/X
+ VGND VGND VPWR VPWR __dut__._1248_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1655__A __dut__.__uuf__._2008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_60_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1127_ __dut__._1129_/A1 __dut__._1127_/A2 __dut__._1126_/X VGND VGND VPWR
+ VPWR __dut__._1127_/X sky130_fd_sc_hd__a21o_4
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1058_ __dut__._1766_/A __dut__._1058_/B VGND VGND VPWR VPWR __dut__._1058_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_98_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_122_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2099__CLK __dut__.__uuf__._2164_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1500_ __dut__.__uuf__._1487_/X __dut__.__uuf__._1483_/X __dut__._1176_/B
+ __dut__.__uuf__._1493_/X __dut__.__uuf__._1499_/X VGND VGND VPWR VPWR __dut__._1175_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1431_ __dut__.__uuf__._1070_/X __dut__.__uuf__._1430_/X __dut__._1206_/B
+ __dut__.__uuf__._1070_/X VGND VGND VPWR VPWR __dut__._1205_/A2 sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._0905__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1362_ __dut__.__uuf__._1367_/A VGND VGND VPWR VPWR __dut__.__uuf__._1362_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1293_ __dut__.__uuf__._1316_/A VGND VGND VPWR VPWR __dut__.__uuf__._1293_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_85_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1633__A2 mc[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1629_ __dut__.__uuf__._1630_/A VGND VGND VPWR VPWR __dut__.__uuf__._1629_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._0922__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1814_ clkbuf_4_6_0_tck/X __dut__._1814_/D __dut__._1515_/Y VGND VGND VPWR
+ VPWR __dut__._1814_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1745_ __dut__._1543_/Y mp[23] __dut__._1744_/X VGND VGND VPWR VPWR __dut__._1745_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1676_ __dut__._1788_/A __dut__._1823_/Q VGND VGND VPWR VPWR __dut__._1676_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1853__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1980_ __dut__.__uuf__._1990_/A __dut__.__uuf__._1980_/B __dut__.__uuf__._1980_/C
+ VGND VGND VPWR VPWR __dut__._1119_/A2 sky130_fd_sc_hd__and3_4
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1379__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1414_ __dut__._1214_/B VGND VGND VPWR VPWR __dut__.__uuf__._1414_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1551__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2114__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1345_ __dut__.__uuf__._1340_/X __dut__.__uuf__._1344_/X __dut__._1240_/B
+ __dut__.__uuf__._1340_/X VGND VGND VPWR VPWR __dut__._1239_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1530_ rst VGND VGND VPWR VPWR __dut__._1530_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1276_ __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR __dut__.__uuf__._1276_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1461_ rst VGND VGND VPWR VPWR __dut__._1461_/Y sky130_fd_sc_hd__inv_2
X__dut__._1392_ __dut__._1542_/A prod[61] VGND VGND VPWR VPWR __dut__._1392_/X sky130_fd_sc_hd__and2_4
XFILLER_46_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1876__CLK __dut__._1919_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpsn_inst_psn_buff_1 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0921_/A1 sky130_fd_sc_hd__buf_2
X_271_ _314_/CLK _271_/D VGND VGND VPWR VPWR _271_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_psn_inst_psn_buff_23_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1748__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1728_ __dut__._1788_/A __dut__._1836_/Q VGND VGND VPWR VPWR __dut__._1728_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1483__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1659_ __dut__._1767_/A1 __dut__._1657_/X __dut__._1658_/X VGND VGND VPWR
+ VPWR __dut__._1818_/D sky130_fd_sc_hd__a21o_4
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1658__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1781__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1130_ __dut__.__uuf__._1130_/A VGND VGND VPWR VPWR __dut__.__uuf__._1130_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1061_ __dut__.__uuf__._1061_/A __dut__.__uuf__._1061_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1061_/Y sky130_fd_sc_hd__nand2_4
XFILLER_83_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1899__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1963_ __dut__._1677_/X VGND VGND VPWR VPWR __dut__.__uuf__._1968_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_36_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1894_ __dut__.__uuf__._1881_/X __dut__.__uuf__._1893_/B __dut__.__uuf__._1893_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1895_/C sky130_fd_sc_hd__o21ai_4
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1568__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_30 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1285_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._0961_ __dut__._0961_/A1 prod[12] __dut__._0960_/X VGND VGND VPWR VPWR __dut__._1897_/D
+ sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_41 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._0991_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_74 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1039_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_63 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1159_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_52 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1771_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._0892_ __dut__._1378_/A __dut__._1862_/Q VGND VGND VPWR VPWR __dut__._0892_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_96 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1116_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_85 psn_inst_psn_buff_88/A VGND VGND VPWR VPWR __dut__._1275_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1328_ __dut__.__uuf__._1328_/A VGND VGND VPWR VPWR __dut__.__uuf__._1380_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1513_ rst VGND VGND VPWR VPWR __dut__._1513_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1259_ __dut__.__uuf__._1263_/A VGND VGND VPWR VPWR __dut__.__uuf__._1259_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_74_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1444_ rst VGND VGND VPWR VPWR __dut__._1444_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1375_ __dut__._1383_/A1 __dut__._1375_/A2 __dut__._1374_/X VGND VGND VPWR
+ VPWR __dut__._1375_/X sky130_fd_sc_hd__a21o_4
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_254_ _199_/A _307_/Q VGND VGND VPWR VPWR _254_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1478__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_185_ _268_/Q _187_/B VGND VGND VPWR VPWR _267_/D sky130_fd_sc_hd__or2_4
XFILLER_89_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1388__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2162_ __dut__.__uuf__._2164_/CLK __dut__._1313_/X __dut__.__uuf__._1200_/X
+ VGND VGND VPWR VPWR prod[22] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1113_ __dut__.__uuf__._1115_/A VGND VGND VPWR VPWR __dut__.__uuf__._1113_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2093_ __dut__.__uuf__._2107_/CLK __dut__._1175_/X __dut__.__uuf__._1498_/X
+ VGND VGND VPWR VPWR __dut__._1176_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1044_ __dut__.__uuf__._1100_/A __dut__.__uuf__._1036_/X __dut__.__uuf__._1037_/X
+ __dut__._0936_/B __dut__.__uuf__._1043_/X VGND VGND VPWR VPWR __dut__._1409_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_68_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1160_ __dut__._1766_/A __dut__._1160_/B VGND VGND VPWR VPWR __dut__._1160_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1946_ __dut__.__uuf__._1946_/A VGND VGND VPWR VPWR __dut__.__uuf__._1990_/A
+ sky130_fd_sc_hd__buf_2
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1091_ __dut__._1129_/A1 __dut__._1091_/A2 __dut__._1090_/X VGND VGND VPWR
+ VPWR __dut__._1091_/X sky130_fd_sc_hd__a21o_4
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1877_ __dut__.__uuf__._1873_/Y __dut__.__uuf__._1874_/Y __dut__.__uuf__._1831_/X
+ __dut__.__uuf__._1876_/X VGND VGND VPWR VPWR __dut__.__uuf__._1878_/A sky130_fd_sc_hd__a211o_4
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1745__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1914__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0944_ __dut__._0944_/A __dut__._1888_/Q VGND VGND VPWR VPWR __dut__._0944_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._0930__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0875_ __dut__._1767_/A1 __dut__._0873_/X __dut__._0874_/X VGND VGND VPWR
+ VPWR __dut__._1854_/D sky130_fd_sc_hd__a21o_4
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_90_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1427_ rst VGND VGND VPWR VPWR __dut__._1427_/Y sky130_fd_sc_hd__inv_2
X__dut__._1358_ __dut__._1378_/A prod[44] VGND VGND VPWR VPWR __dut__._1358_/X sky130_fd_sc_hd__and2_4
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1289_ __dut__._1289_/A1 __dut__._1289_/A2 __dut__._1288_/X VGND VGND VPWR
+ VPWR __dut__._1289_/X sky130_fd_sc_hd__a21o_4
XFILLER_91_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_306_ _306_/CLK _306_/D trst VGND VGND VPWR VPWR _306_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_237_ _237_/A _313_/Q VGND VGND VPWR VPWR _238_/D sky130_fd_sc_hd__nor2_4
X_168_ _282_/Q _173_/B VGND VGND VPWR VPWR _281_/D sky130_fd_sc_hd__and2_4
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_152_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1390__B prod[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1800_ __dut__.__uuf__._1796_/Y __dut__.__uuf__._1797_/Y __dut__.__uuf__._1798_/X
+ __dut__.__uuf__._1804_/B VGND VGND VPWR VPWR __dut__.__uuf__._1800_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1731_ __dut__._1034_/B VGND VGND VPWR VPWR __dut__.__uuf__._1731_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1662_ __dut__._1637_/X VGND VGND VPWR VPWR __dut__.__uuf__._1670_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1593_ __dut__.__uuf__._1593_/A VGND VGND VPWR VPWR __dut__.__uuf__._1593_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2145_ __dut__.__uuf__._2164_/CLK __dut__._1279_/X __dut__.__uuf__._1248_/X
+ VGND VGND VPWR VPWR prod[5] sky130_fd_sc_hd__dfrtp_4
XFILLER_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2076_ __dut__.__uuf__._2107_/CLK __dut__._1141_/X __dut__.__uuf__._1565_/X
+ VGND VGND VPWR VPWR __dut__._1142_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1027_ __dut__._1402_/B VGND VGND VPWR VPWR __dut__.__uuf__._1061_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1212_ __dut__._1786_/A __dut__._1212_/B VGND VGND VPWR VPWR __dut__._1212_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1143_ __dut__._1647_/A1 __dut__._1143_/A2 __dut__._1142_/X VGND VGND VPWR
+ VPWR __dut__._1143_/X sky130_fd_sc_hd__a21o_4
XANTENNA__286__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1929_ __dut__._1100_/B VGND VGND VPWR VPWR __dut__.__uuf__._1929_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1074_ __dut__._1074_/A __dut__._1074_/B VGND VGND VPWR VPWR __dut__._1074_/X
+ sky130_fd_sc_hd__and2_4
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._0927_ __dut__._1395_/A1 prod[60] __dut__._0926_/X VGND VGND VPWR VPWR __dut__._1880_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1756__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._0941__A2 prod[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__299__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1491__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1709__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1666__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1714_ __dut__.__uuf__._1908_/A VGND VGND VPWR VPWR __dut__.__uuf__._1936_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_21_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1645_ __dut__.__uuf__._1648_/A VGND VGND VPWR VPWR __dut__.__uuf__._1645_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1830_ clkbuf_4_7_0_tck/X __dut__._1830_/D __dut__._1499_/Y VGND VGND VPWR
+ VPWR __dut__._1830_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1576_ __dut__.__uuf__._1580_/A VGND VGND VPWR VPWR __dut__.__uuf__._1576_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1576__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1761_ __dut__._1543_/Y mp[27] __dut__._1760_/X VGND VGND VPWR VPWR __dut__._1761_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1692_ __dut__._1788_/A __dut__._1827_/Q VGND VGND VPWR VPWR __dut__._1692_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2128_ __dut__.__uuf__._2206_/CLK __dut__._1245_/X __dut__.__uuf__._1327_/X
+ VGND VGND VPWR VPWR __dut__._1246_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2059_ __dut__.__uuf__._2065_/CLK __dut__._1107_/X __dut__.__uuf__._1595_/X
+ VGND VGND VPWR VPWR __dut__._1108_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_53_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1126_ __dut__._1678_/A __dut__._1126_/B VGND VGND VPWR VPWR __dut__._1126_/X
+ sky130_fd_sc_hd__and2_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1057_ __dut__._1057_/A1 __dut__._1057_/A2 __dut__._1056_/X VGND VGND VPWR
+ VPWR __dut__._1057_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2020__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1486__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__301__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_115_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1581__A __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1430_ __dut__.__uuf__._1429_/Y __dut__.__uuf__._1425_/X __dut__.__uuf__._1324_/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._1430_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1361_ __dut__.__uuf__._1354_/X __dut__.__uuf__._1360_/X __dut__._1234_/B
+ __dut__.__uuf__._1354_/X VGND VGND VPWR VPWR __dut__._1233_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1292_ __dut__.__uuf__._1346_/A VGND VGND VPWR VPWR __dut__.__uuf__._1316_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_tck clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR clkbuf_3_7_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1628_ __dut__.__uuf__._1630_/A VGND VGND VPWR VPWR __dut__.__uuf__._1628_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1813_ clkbuf_4_6_0_tck/X __dut__._1813_/D __dut__._1516_/Y VGND VGND VPWR
+ VPWR __dut__._1813_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1559_ __dut__.__uuf__._1569_/A VGND VGND VPWR VPWR __dut__.__uuf__._1559_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1744_ __dut__._1788_/A __dut__._1840_/Q VGND VGND VPWR VPWR __dut__._1744_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1675_ __dut__._1767_/A1 __dut__._1673_/X __dut__._1674_/X VGND VGND VPWR
+ VPWR __dut__._1822_/D sky130_fd_sc_hd__a21o_4
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1085__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0___dut__.__uuf__.__clk_source__ clkbuf_4_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2083_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__._1109_ __dut__._1129_/A1 __dut__._1109_/A2 __dut__._1108_/X VGND VGND VPWR
+ VPWR __dut__._1109_/X sky130_fd_sc_hd__a21o_4
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0899__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2066__CLK __dut__.__uuf__._2119_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1413_ __dut__.__uuf__._1418_/A VGND VGND VPWR VPWR __dut__.__uuf__._1413_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1344_ __dut__.__uuf__._1343_/Y __dut__.__uuf__._1323_/X __dut__.__uuf__._1324_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1344_/X sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._1551__A2 __dut__._1549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1275_ __dut__.__uuf__._1295_/A VGND VGND VPWR VPWR __dut__.__uuf__._1495_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_100_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1460_ rst VGND VGND VPWR VPWR __dut__._1460_/Y sky130_fd_sc_hd__inv_2
X__dut__._1391_ __dut__._1395_/A1 __dut__._1391_/A2 __dut__._1390_/X VGND VGND VPWR
+ VPWR __dut__._1391_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_2 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1383_/A1 sky130_fd_sc_hd__buf_8
XANTENNA__255__D tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_270_ _314_/CLK _270_/D VGND VGND VPWR VPWR _270_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_psn_inst_psn_buff_16_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1764__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1727_ __dut__._1727_/A1 __dut__._1725_/X __dut__._1726_/X VGND VGND VPWR
+ VPWR __dut__._1835_/D sky130_fd_sc_hd__a21o_4
X__dut__._1658_ __dut__._1766_/A __dut__._1817_/Q VGND VGND VPWR VPWR __dut__._1658_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1589_ __dut__._1543_/Y mc[1] __dut__._1588_/X VGND VGND VPWR VPWR __dut__._1589_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_17_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1781__A2 mp[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1674__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1060_ __dut__.__uuf__._1063_/A VGND VGND VPWR VPWR __dut__.__uuf__._1060_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1962_ __dut__._1112_/B VGND VGND VPWR VPWR __dut__.__uuf__._1962_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1893_ __dut__.__uuf__._1914_/A __dut__.__uuf__._1893_/B __dut__.__uuf__._1893_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1895_/B sky130_fd_sc_hd__or3_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1221__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_31 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR psn_inst_psn_buff_49/A
+ sky130_fd_sc_hd__buf_8
X__dut__._0960_ __dut__._1324_/A __dut__._1896_/Q VGND VGND VPWR VPWR __dut__._0960_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_20 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0939_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_42 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._0993_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_64 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1153_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_53 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1763_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__._0891_ __dut__._1383_/A1 prod[42] __dut__._0890_/X VGND VGND VPWR VPWR __dut__._1862_/D
+ sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_75 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1037_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_97 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1112_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_86 psn_inst_psn_buff_88/A VGND VGND VPWR VPWR __dut__._1197_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1327_ __dut__.__uuf__._1342_/A VGND VGND VPWR VPWR __dut__.__uuf__._1327_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1584__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1512_ rst VGND VGND VPWR VPWR __dut__._1512_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1258_ __dut__.__uuf__._1257_/X __dut__.__uuf__._1254_/X prod[3]
+ prod[4] __dut__.__uuf__._1249_/X VGND VGND VPWR VPWR __dut__._1275_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1189_ __dut__.__uuf__._1189_/A VGND VGND VPWR VPWR __dut__.__uuf__._1189_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1443_ rst VGND VGND VPWR VPWR __dut__._1443_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1843__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1374_ __dut__._1378_/A prod[52] VGND VGND VPWR VPWR __dut__._1374_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._0928__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_253_ _196_/X _259_/Q VGND VGND VPWR VPWR _253_/Q sky130_fd_sc_hd__dfxtp_4
X_184_ _269_/Q _191_/B VGND VGND VPWR VPWR _268_/D sky130_fd_sc_hd__and2_4
XFILLER_89_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1494__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2104__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1388__B prod[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2161_ __dut__.__uuf__._2210_/CLK __dut__._1311_/X __dut__.__uuf__._1202_/X
+ VGND VGND VPWR VPWR prod[21] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1112_ __dut__.__uuf__._1109_/X __dut__.__uuf__._1106_/X prod[52]
+ prod[53] __dut__.__uuf__._1100_/X VGND VGND VPWR VPWR __dut__._1373_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1866__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2092_ __dut__.__uuf__._2107_/CLK __dut__._1173_/X __dut__.__uuf__._1501_/X
+ VGND VGND VPWR VPWR __dut__._1174_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1043_ __dut__.__uuf__._1416_/A VGND VGND VPWR VPWR __dut__.__uuf__._1043_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1090_ __dut__._1094_/A __dut__._1090_/B VGND VGND VPWR VPWR __dut__._1090_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1945_ __dut__.__uuf__._1945_/A VGND VGND VPWR VPWR __dut__._1109_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1876_ __dut__.__uuf__._1873_/Y __dut__.__uuf__._1874_/Y __dut__.__uuf__._1853_/X
+ __dut__.__uuf__._1880_/B VGND VGND VPWR VPWR __dut__.__uuf__._1876_/X sky130_fd_sc_hd__o22a_4
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1745__A2 mp[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0943_ __dut__._0943_/A1 prod[3] __dut__._0942_/X VGND VGND VPWR VPWR __dut__._1888_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0874_ __dut__._1766_/A __dut__._1853_/Q VGND VGND VPWR VPWR __dut__._0874_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_78_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_83_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1681__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1426_ rst VGND VGND VPWR VPWR __dut__._1426_/Y sky130_fd_sc_hd__inv_2
X__dut__._1357_ __dut__._1383_/A1 __dut__._1357_/A2 __dut__._1356_/X VGND VGND VPWR
+ VPWR __dut__._1357_/X sky130_fd_sc_hd__a21o_4
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1288_ __dut__._1770_/A prod[9] VGND VGND VPWR VPWR __dut__._1288_/X sky130_fd_sc_hd__and2_4
XFILLER_91_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_305_ _306_/CLK _305_/D trst VGND VGND VPWR VPWR _305_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1489__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_236_ _305_/Q _306_/Q VGND VGND VPWR VPWR _236_/Y sky130_fd_sc_hd__nor2_4
X_167_ _283_/Q _172_/B VGND VGND VPWR VPWR _282_/D sky130_fd_sc_hd__or2_4
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1889__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_145_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1730_ __dut__.__uuf__._1773_/A __dut__.__uuf__._1730_/B __dut__.__uuf__._1730_/C
+ VGND VGND VPWR VPWR __dut__._1027_/A2 sky130_fd_sc_hd__and3_4
X__dut__.__uuf__._1661_ __dut__.__uuf__._1908_/A VGND VGND VPWR VPWR __dut__.__uuf__._2001_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1592_ __dut__.__uuf__._1593_/A VGND VGND VPWR VPWR __dut__.__uuf__._1592_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2144_ __dut__.__uuf__._2208_/CLK __dut__._1277_/X __dut__.__uuf__._1253_/X
+ VGND VGND VPWR VPWR prod[4] sky130_fd_sc_hd__dfrtp_4
XFILLER_75_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2075_ __dut__.__uuf__._2107_/CLK __dut__._1139_/X __dut__.__uuf__._1569_/X
+ VGND VGND VPWR VPWR __dut__._1140_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1494__A __dut__.__uuf__._1536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1026_ __dut__.__uuf__._1190_/A VGND VGND VPWR VPWR __dut__.__uuf__._1100_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1663__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1211_ __dut__._1787_/A1 __dut__._1211_/A2 __dut__._1210_/X VGND VGND VPWR
+ VPWR __dut__._1211_/X sky130_fd_sc_hd__a21o_4
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1142_ __dut__._1142_/A __dut__._1142_/B VGND VGND VPWR VPWR __dut__._1142_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1928_ __dut__._1106_/B VGND VGND VPWR VPWR __dut__.__uuf__._1928_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1073_ __dut__._1129_/A1 __dut__._1073_/A2 __dut__._1072_/X VGND VGND VPWR
+ VPWR __dut__._1073_/X sky130_fd_sc_hd__a21o_4
XFILLER_51_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1859_ __dut__.__uuf__._1859_/A __dut__.__uuf__._1859_/B __dut__.__uuf__._1859_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1861_/B sky130_fd_sc_hd__or3_4
XFILLER_8_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._0926_ __dut__._1542_/A __dut__._1879_/Q VGND VGND VPWR VPWR __dut__._0926_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1772__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1409_ __dut__._1409_/A1 __dut__._1409_/A2 __dut__._1408_/X VGND VGND VPWR
+ VPWR __dut__._1409_/X sky130_fd_sc_hd__a21o_4
XFILLER_74_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1709__A2 mp[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ _294_/Q _293_/Q _222_/A VGND VGND VPWR VPWR _293_/D sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._1682__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1645__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1713_ __dut__.__uuf__._1749_/A __dut__.__uuf__._1713_/B __dut__.__uuf__._1713_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1717_/B sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1644_ __dut__.__uuf__._1648_/A VGND VGND VPWR VPWR __dut__.__uuf__._1644_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1575_ __dut__.__uuf__._1575_/A VGND VGND VPWR VPWR __dut__.__uuf__._1580_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1760_ __dut__._1788_/A __dut__._1844_/Q VGND VGND VPWR VPWR __dut__._1760_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1691_ __dut__._1719_/A1 __dut__._1689_/X __dut__._1690_/X VGND VGND VPWR
+ VPWR __dut__._1826_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._2127_ __dut__.__uuf__._2206_/CLK __dut__._1243_/X __dut__.__uuf__._1333_/X
+ VGND VGND VPWR VPWR __dut__._1244_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1592__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2058_ __dut__.__uuf__._2065_/CLK __dut__._1105_/X __dut__.__uuf__._1596_/X
+ VGND VGND VPWR VPWR __dut__._1106_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_tck tck VGND VGND VPWR VPWR clkbuf_0_tck/X sky130_fd_sc_hd__clkbuf_16
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_46_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1125_ __dut__._1129_/A1 __dut__._1125_/A2 __dut__._1124_/X VGND VGND VPWR
+ VPWR __dut__._1125_/X sky130_fd_sc_hd__a21o_4
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1056_ __dut__._1056_/A __dut__._1056_/B VGND VGND VPWR VPWR __dut__._1056_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._0909_ __dut__._1383_/A1 prod[51] __dut__._0908_/X VGND VGND VPWR VPWR __dut__._1871_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1889_ __dut__._1902_/CLK __dut__._1889_/D __dut__._1440_/Y VGND VGND VPWR
+ VPWR __dut__._1889_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1627__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_108_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1396__B prod[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1360_ __dut__.__uuf__._1359_/Y __dut__.__uuf__._1349_/X __dut__.__uuf__._1350_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1360_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1291_ __dut__.__uuf__._1286_/X __dut__.__uuf__._1290_/X __dut__._1260_/B
+ __dut__.__uuf__._1286_/X VGND VGND VPWR VPWR __dut__._1259_/A2 sky130_fd_sc_hd__a2bb2o_4
XANTENNA__276__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1627_ __dut__.__uuf__._1630_/A VGND VGND VPWR VPWR __dut__.__uuf__._1627_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1812_ clkbuf_4_6_0_tck/X __dut__._1812_/D __dut__._1517_/Y VGND VGND VPWR
+ VPWR __dut__._1812_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1558_ __dut__.__uuf__._1551_/X __dut__.__uuf__._1547_/X __dut__._1148_/B
+ __dut__.__uuf__._1449_/A __dut__.__uuf__._1557_/X VGND VGND VPWR VPWR __dut__._1147_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1489_ __dut__.__uuf__._1487_/X __dut__.__uuf__._1483_/X __dut__._1180_/B
+ __dut__.__uuf__._1471_/X __dut__.__uuf__._1488_/X VGND VGND VPWR VPWR __dut__._1179_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1743_ __dut__._1759_/A1 __dut__._1741_/X __dut__._1742_/X VGND VGND VPWR
+ VPWR __dut__._1839_/D sky130_fd_sc_hd__a21o_4
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1674_ __dut__._1766_/A __dut__._1821_/Q VGND VGND VPWR VPWR __dut__._1674_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1609__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1444__A2 __dut__.__uuf__._1946_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1108_ __dut__._1108_/A __dut__._1108_/B VGND VGND VPWR VPWR __dut__._1108_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1039_ __dut__._1039_/A1 __dut__._1039_/A2 __dut__._1038_/X VGND VGND VPWR
+ VPWR __dut__._1039_/X sky130_fd_sc_hd__a21o_4
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1497__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__299__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1412_ __dut__.__uuf__._1405_/X __dut__.__uuf__._1411_/X __dut__._1214_/B
+ __dut__.__uuf__._1405_/X VGND VGND VPWR VPWR __dut__._1213_/A2 sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_4_15_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2194_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1343_ __dut__._1242_/B VGND VGND VPWR VPWR __dut__.__uuf__._1343_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1274_ __dut__.__uuf__._1314_/A VGND VGND VPWR VPWR __dut__.__uuf__._1274_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1390_ __dut__._1542_/A prod[60] VGND VGND VPWR VPWR __dut__._1390_/X sky130_fd_sc_hd__and2_4
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2010__CLK __dut__.__uuf__._2119_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2160__CLK __dut__.__uuf__._2164_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_14_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_3 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1385_/A1 sky130_fd_sc_hd__buf_2
XFILLER_22_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1110__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1726_ __dut__._1766_/A __dut__._1833_/Q VGND VGND VPWR VPWR __dut__._1726_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_89_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1657_ __dut__._1543_/Y mp[3] __dut__._1656_/X VGND VGND VPWR VPWR __dut__._1657_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1588_ __dut__._1788_/A __dut__._1801_/Q VGND VGND VPWR VPWR __dut__._1588_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1780__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_tck clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR clkbuf_3_5_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2033__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1690__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__314__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1961_ __dut__._1118_/B VGND VGND VPWR VPWR __dut__.__uuf__._1961_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1892_ __dut__.__uuf__._1884_/Y __dut__.__uuf__._1885_/Y __dut__.__uuf__._1884_/Y
+ __dut__.__uuf__._1885_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1893_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._1795__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_10 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1341_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_21 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1787_/A1
+ sky130_fd_sc_hd__buf_8
X__dut__._0890_ __dut__._1378_/A __dut__._1861_/Q VGND VGND VPWR VPWR __dut__._0890_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_43 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._1325_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_65 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1155_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_54 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1739_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_32 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._0951_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_98 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1108_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_76 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1075_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_87 psn_inst_psn_buff_88/A VGND VGND VPWR VPWR __dut__._1193_/A1
+ sky130_fd_sc_hd__buf_8
X__dut__.__uuf__._1326_ __dut__.__uuf__._1314_/X __dut__.__uuf__._1325_/X __dut__._1248_/B
+ __dut__.__uuf__._1314_/X VGND VGND VPWR VPWR __dut__._1247_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1511_ rst VGND VGND VPWR VPWR __dut__._1511_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1257_ __dut__.__uuf__._1466_/A VGND VGND VPWR VPWR __dut__.__uuf__._1257_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1188_ __dut__.__uuf__._1183_/X __dut__.__uuf__._1180_/X prod[26]
+ prod[27] __dut__.__uuf__._1175_/X VGND VGND VPWR VPWR __dut__._1321_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1442_ rst VGND VGND VPWR VPWR __dut__._1442_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1373_ __dut__._1383_/A1 __dut__._1373_/A2 __dut__._1372_/X VGND VGND VPWR
+ VPWR __dut__._1373_/X sky130_fd_sc_hd__a21o_4
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_252_ _197_/X _315_/Q VGND VGND VPWR VPWR _252_/Q sky130_fd_sc_hd__dfxtp_4
X_183_ _183_/A VGND VGND VPWR VPWR _191_/B sky130_fd_sc_hd__buf_2
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1709_ __dut__._1543_/Y mp[15] __dut__._1708_/X VGND VGND VPWR VPWR __dut__._1709_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1574__B2 __dut__.__uuf__._1069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2160_ __dut__.__uuf__._2164_/CLK __dut__._1309_/X __dut__.__uuf__._1204_/X
+ VGND VGND VPWR VPWR prod[20] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1111_ __dut__.__uuf__._1115_/A VGND VGND VPWR VPWR __dut__.__uuf__._1111_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2091_ __dut__.__uuf__._2107_/CLK __dut__._1171_/X __dut__.__uuf__._1504_/X
+ VGND VGND VPWR VPWR __dut__._1172_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1042_ __dut__.__uuf__._1328_/A VGND VGND VPWR VPWR __dut__.__uuf__._1416_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1944_ __dut__.__uuf__._1939_/Y __dut__.__uuf__._1940_/Y __dut__.__uuf__._1941_/X
+ __dut__.__uuf__._1943_/X VGND VGND VPWR VPWR __dut__.__uuf__._1945_/A sky130_fd_sc_hd__a211o_4
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1875_ __dut__._1553_/X VGND VGND VPWR VPWR __dut__.__uuf__._1880_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2079__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1262__B1 prod[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0942_ __dut__._0942_/A __dut__._1887_/Q VGND VGND VPWR VPWR __dut__._0942_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._0873_ __dut__._1543_/Y mc[9] __dut__._0872_/X VGND VGND VPWR VPWR __dut__._0873_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA__315__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1309_ __dut__.__uuf__._1308_/Y __dut__.__uuf__._1297_/X __dut__.__uuf__._1299_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1309_/X sky130_fd_sc_hd__o21a_4
XANTENNA_psn_inst_psn_buff_76_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1681__A2 mp[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1425_ rst VGND VGND VPWR VPWR __dut__._1425_/Y sky130_fd_sc_hd__inv_2
X__dut__._1356_ __dut__._1378_/A prod[43] VGND VGND VPWR VPWR __dut__._1356_/X sky130_fd_sc_hd__and2_4
X__dut__._1287_ __dut__._1289_/A1 __dut__._1287_/A2 __dut__._1286_/X VGND VGND VPWR
+ VPWR __dut__._1287_/X sky130_fd_sc_hd__a21o_4
X_304_ _306_/CLK _304_/D trst VGND VGND VPWR VPWR _304_/Q sky130_fd_sc_hd__dfrtp_4
X_235_ _251_/Q VGND VGND VPWR VPWR tdo_paden_o sky130_fd_sc_hd__inv_2
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_166_ _284_/Q _173_/B VGND VGND VPWR VPWR _283_/D sky130_fd_sc_hd__and2_4
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1121__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_138_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1660_ __dut__.__uuf__._1660_/A VGND VGND VPWR VPWR __dut__.__uuf__._1660_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1591_ __dut__.__uuf__._1593_/A VGND VGND VPWR VPWR __dut__.__uuf__._1591_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2143_ __dut__.__uuf__._2208_/CLK __dut__._1275_/X __dut__.__uuf__._1256_/X
+ VGND VGND VPWR VPWR prod[3] sky130_fd_sc_hd__dfrtp_4
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2074_ __dut__.__uuf__._2107_/CLK __dut__._1137_/X __dut__.__uuf__._1576_/X
+ VGND VGND VPWR VPWR __dut__._1138_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1025_ __dut__.__uuf__._1226_/A VGND VGND VPWR VPWR __dut__.__uuf__._1190_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1210_ __dut__._1786_/A __dut__._1210_/B VGND VGND VPWR VPWR __dut__._1210_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1141_ __dut__._1647_/A1 __dut__._1141_/A2 __dut__._1140_/X VGND VGND VPWR
+ VPWR __dut__._1141_/X sky130_fd_sc_hd__a21o_4
XFILLER_45_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1927_ __dut__.__uuf__._1938_/A __dut__.__uuf__._1927_/B __dut__.__uuf__._1927_/C
+ VGND VGND VPWR VPWR __dut__._1099_/A2 sky130_fd_sc_hd__and3_4
X__dut__._1072_ __dut__._1074_/A __dut__._1072_/B VGND VGND VPWR VPWR __dut__._1072_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_101_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1858_ __dut__.__uuf__._1851_/Y __dut__.__uuf__._1852_/Y __dut__.__uuf__._1851_/Y
+ __dut__.__uuf__._1852_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1859_/C sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1789_ __dut__.__uuf__._1786_/Y __dut__.__uuf__._1787_/Y __dut__.__uuf__._1743_/X
+ __dut__.__uuf__._1793_/B VGND VGND VPWR VPWR __dut__.__uuf__._1789_/X sky130_fd_sc_hd__o22a_4
X__dut__._0925_ __dut__._1395_/A1 prod[59] __dut__._0924_/X VGND VGND VPWR VPWR __dut__._1879_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1351__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1103__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1408_ __dut__._1408_/A __dut__._1408_/B VGND VGND VPWR VPWR __dut__._1408_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_47_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1339_ __dut__._1339_/A1 __dut__._1339_/A2 __dut__._1338_/X VGND VGND VPWR
+ VPWR __dut__._1339_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1856__CLK __dut__._1919_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._0917__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_218_ _234_/A VGND VGND VPWR VPWR _222_/A sky130_fd_sc_hd__buf_2
X_149_ _239_/A _142_/Y _309_/Q _308_/Q _144_/Y VGND VGND VPWR VPWR _308_/D sky130_fd_sc_hd__a32o_4
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1645__A2 mp[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1712_ __dut__.__uuf__._1706_/Y __dut__.__uuf__._1707_/Y __dut__.__uuf__._1706_/Y
+ __dut__.__uuf__._1707_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1713_/C sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1643_ __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR __dut__.__uuf__._1648_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1574_ __dut__.__uuf__._1573_/X __dut__.__uuf__._2004_/B __dut__._1142_/B
+ __dut__.__uuf__._1069_/X VGND VGND VPWR VPWR __dut__._1139_/A2 sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._1581__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2117__CLK __dut__.__uuf__._2119_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_88_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1690_ __dut__._1766_/A __dut__._1825_/Q VGND VGND VPWR VPWR __dut__._1690_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2126_ __dut__.__uuf__._2138_/CLK __dut__._1241_/X __dut__.__uuf__._1337_/X
+ VGND VGND VPWR VPWR __dut__._1242_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2057_ __dut__.__uuf__._2065_/CLK __dut__._1103_/X __dut__.__uuf__._1597_/X
+ VGND VGND VPWR VPWR __dut__._1104_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1879__CLK __dut__._1919_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1124_ __dut__._1128_/A __dut__._1124_/B VGND VGND VPWR VPWR __dut__._1124_/X
+ sky130_fd_sc_hd__and2_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_39_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1055_ __dut__._1055_/A1 __dut__._1055_/A2 __dut__._1054_/X VGND VGND VPWR
+ VPWR __dut__._1055_/X sky130_fd_sc_hd__a21o_4
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._0952__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0908_ __dut__._1378_/A __dut__._1870_/Q VGND VGND VPWR VPWR __dut__._0908_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1888_ __dut__._1902_/CLK __dut__._1888_/D __dut__._1441_/Y VGND VGND VPWR
+ VPWR __dut__._1888_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0862__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1563__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1290_ __dut__.__uuf__._1289_/Y __dut__.__uuf__._1276_/X __dut__.__uuf__._1271_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1290_/X sky130_fd_sc_hd__o21a_4
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1626_ __dut__.__uuf__._1630_/A VGND VGND VPWR VPWR __dut__.__uuf__._1626_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1811_ clkbuf_4_6_0_tck/X __dut__._1811_/D __dut__._1518_/Y VGND VGND VPWR
+ VPWR __dut__._1811_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1557_ __dut__._1657_/X __dut__.__uuf__._1078_/A __dut__._1150_/B
+ __dut__.__uuf__._1660_/A VGND VGND VPWR VPWR __dut__.__uuf__._1557_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1488_ __dut__._1729_/X __dut__.__uuf__._1472_/X __dut__._1182_/B
+ __dut__.__uuf__._1473_/X VGND VGND VPWR VPWR __dut__.__uuf__._1488_/X sky130_fd_sc_hd__o22a_4
X__dut__._1742_ __dut__._1770_/A __dut__._1838_/Q VGND VGND VPWR VPWR __dut__._1742_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1673_ __dut__._1543_/Y mp[7] __dut__._1672_/X VGND VGND VPWR VPWR __dut__._1673_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2109_ __dut__.__uuf__._2114_/CLK __dut__._1207_/X __dut__.__uuf__._1423_/X
+ VGND VGND VPWR VPWR __dut__._1208_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_91_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1609__A2 mc[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1107_ __dut__._1129_/A1 __dut__._1107_/A2 __dut__._1106_/X VGND VGND VPWR
+ VPWR __dut__._1107_/X sky130_fd_sc_hd__a21o_4
X__dut__._1038_ __dut__._1678_/A __dut__._1038_/B VGND VGND VPWR VPWR __dut__._1038_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1778__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1545__A1 mc[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_120_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1688__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1411_ __dut__.__uuf__._1410_/Y __dut__.__uuf__._1400_/X __dut__.__uuf__._1401_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1411_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_3_7_0___dut__.__uuf__.__clk_source__ clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0___dut__.__uuf__.__clk_source__/X sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1342_ __dut__.__uuf__._1342_/A VGND VGND VPWR VPWR __dut__.__uuf__._1342_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1273_ __dut__.__uuf__._1288_/A VGND VGND VPWR VPWR __dut__.__uuf__._1273_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpsn_inst_psn_buff_4 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1387_/A1 sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1917__CLK __dut__._1917_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1598__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1609_ __dut__.__uuf__._1611_/A VGND VGND VPWR VPWR __dut__.__uuf__._1609_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_78_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1725_ __dut__._1543_/Y mp[18] __dut__._1724_/X VGND VGND VPWR VPWR __dut__._1725_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1656_ __dut__._1788_/A __dut__._1818_/Q VGND VGND VPWR VPWR __dut__._1656_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1587_ __dut__._1767_/A1 __dut__._1585_/X __dut__._1586_/X VGND VGND VPWR
+ VPWR __dut__._1800_/D sky130_fd_sc_hd__a21o_4
XFILLER_76_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__266__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1050__A1 __dut__.__uuf__._1100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_168_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1960_ __dut__.__uuf__._1990_/A __dut__.__uuf__._1960_/B __dut__.__uuf__._1960_/C
+ VGND VGND VPWR VPWR __dut__._1111_/A2 sky130_fd_sc_hd__and3_4
XFILLER_48_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1891_ __dut__.__uuf__._1946_/A VGND VGND VPWR VPWR __dut__.__uuf__._1938_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1757__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_11 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1005_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_22 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0941_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_44 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._1327_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_55 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1759_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_33 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._0953_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_99 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1106_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_77 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1071_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_66 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1655_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_88 psn_inst_psn_buff_88/A VGND VGND VPWR VPWR __dut__._1779_/A1
+ sky130_fd_sc_hd__buf_8
X__dut__.__uuf__._1325_ __dut__.__uuf__._1322_/Y __dut__.__uuf__._1323_/X __dut__.__uuf__._1324_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1325_/X sky130_fd_sc_hd__o21a_4
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1510_ rst VGND VGND VPWR VPWR __dut__._1510_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1256_ __dut__.__uuf__._1263_/A VGND VGND VPWR VPWR __dut__.__uuf__._1256_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1187_ __dut__.__uuf__._1189_/A VGND VGND VPWR VPWR __dut__.__uuf__._1187_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1441_ rst VGND VGND VPWR VPWR __dut__._1441_/Y sky130_fd_sc_hd__inv_2
X__dut__._1372_ __dut__._1378_/A prod[51] VGND VGND VPWR VPWR __dut__._1372_/X sky130_fd_sc_hd__and2_4
XFILLER_39_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__289__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_251_ _198_/X _251_/D VGND VGND VPWR VPWR _251_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_21_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_182_ _270_/Q _182_/B VGND VGND VPWR VPWR _269_/D sky130_fd_sc_hd__and2_4
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1708_ __dut__._1788_/A __dut__._1831_/Q VGND VGND VPWR VPWR __dut__._1708_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1639_ __dut__._1647_/A1 __dut__._1637_/X __dut__._1638_/X VGND VGND VPWR
+ VPWR __dut__._1813_/D sky130_fd_sc_hd__a21o_4
XFILLER_18_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._0870__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1110_ __dut__.__uuf__._1109_/X __dut__.__uuf__._1106_/X prod[53]
+ prod[54] __dut__.__uuf__._1100_/X VGND VGND VPWR VPWR __dut__._1375_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2090_ __dut__.__uuf__._2097_/CLK __dut__._1169_/X __dut__.__uuf__._1508_/X
+ VGND VGND VPWR VPWR __dut__._1170_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1041_ __dut__.__uuf__._1448_/A VGND VGND VPWR VPWR __dut__.__uuf__._1328_/A
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1206__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1943_ __dut__.__uuf__._1939_/Y __dut__.__uuf__._1940_/Y __dut__.__uuf__._1908_/X
+ __dut__.__uuf__._1948_/B VGND VGND VPWR VPWR __dut__.__uuf__._1943_/X sky130_fd_sc_hd__o22a_4
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1874_ __dut__._1080_/B VGND VGND VPWR VPWR __dut__.__uuf__._1874_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._0941_ __dut__._0941_/A1 prod[2] __dut__._0940_/X VGND VGND VPWR VPWR __dut__._1887_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0872_ __dut__._1788_/A __dut__._1854_/Q VGND VGND VPWR VPWR __dut__._0872_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1308_ __dut__._1256_/B VGND VGND VPWR VPWR __dut__.__uuf__._1308_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1239_ __dut__.__uuf__._1483_/A VGND VGND VPWR VPWR __dut__.__uuf__._1239_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1424_ rst VGND VGND VPWR VPWR __dut__._1424_/Y sky130_fd_sc_hd__inv_2
X__dut__._1355_ __dut__._1383_/A1 __dut__._1355_/A2 __dut__._1354_/X VGND VGND VPWR
+ VPWR __dut__._1355_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_69_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_tck clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR clkbuf_3_3_0_tck/A sky130_fd_sc_hd__clkbuf_1
X__dut__._1286_ __dut__._1770_/A prod[8] VGND VGND VPWR VPWR __dut__._1286_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2023__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_303_ _306_/CLK _303_/D trst VGND VGND VPWR VPWR _303_/Q sky130_fd_sc_hd__dfrtp_4
X_234_ _234_/A _234_/B VGND VGND VPWR VPWR _305_/D sky130_fd_sc_hd__and2_4
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1786__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_165_ _183_/A VGND VGND VPWR VPWR _173_/B sky130_fd_sc_hd__buf_2
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1590_ __dut__.__uuf__._1593_/A VGND VGND VPWR VPWR __dut__.__uuf__._1590_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._0935__A2 done VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1696__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2142_ __dut__.__uuf__._2208_/CLK __dut__._1273_/X __dut__.__uuf__._1259_/X
+ VGND VGND VPWR VPWR prod[2] sky130_fd_sc_hd__dfrtp_4
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2073_ __dut__.__uuf__._2107_/CLK __dut__._1135_/X __dut__.__uuf__._1577_/X
+ VGND VGND VPWR VPWR __dut__._1136_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1024_ __dut__.__uuf__._2005_/A __dut__._1138_/B __dut__.__uuf__._1024_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1226_/A sky130_fd_sc_hd__or3_4
XFILLER_83_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0871__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2046__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1140_ __dut__._1140_/A __dut__._1140_/B VGND VGND VPWR VPWR __dut__._1140_/X
+ sky130_fd_sc_hd__and2_4
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1926_ __dut__.__uuf__._1881_/X __dut__.__uuf__._1925_/B __dut__.__uuf__._1925_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1927_/C sky130_fd_sc_hd__o21ai_4
X__dut__._1071_ __dut__._1071_/A1 __dut__._1071_/A2 __dut__._1070_/X VGND VGND VPWR
+ VPWR __dut__._1071_/X sky130_fd_sc_hd__a21o_4
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1857_ __dut__.__uuf__._1857_/A VGND VGND VPWR VPWR __dut__._1077_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_61_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1788_ __dut__._1585_/X VGND VGND VPWR VPWR __dut__.__uuf__._1793_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._0924_ __dut__._1542_/A __dut__._1878_/Q VGND VGND VPWR VPWR __dut__._0924_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1407_ __dut__._1409_/A1 __dut__._1407_/A2 __dut__._1406_/X VGND VGND VPWR
+ VPWR __dut__._1407_/X sky130_fd_sc_hd__a21o_4
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1338_ __dut__._1338_/A prod[34] VGND VGND VPWR VPWR __dut__._1338_/X sky130_fd_sc_hd__and2_4
X__dut__._1269_ __dut__._1787_/A1 __dut__._1269_/A2 __dut__._1268_/X VGND VGND VPWR
+ VPWR __dut__._1269_/X sky130_fd_sc_hd__a21o_4
XFILLER_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_217_ _293_/Q _232_/A VGND VGND VPWR VPWR _292_/D sky130_fd_sc_hd__and2_4
X_148_ _309_/Q _146_/Y _296_/Q _147_/X VGND VGND VPWR VPWR _309_/D sky130_fd_sc_hd__a211o_4
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_150_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2069__CLK __dut__.__uuf__._2119_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_65_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1800__CLK __dut__._1410_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1711_ __dut__.__uuf__._1711_/A VGND VGND VPWR VPWR __dut__._1025_/A2
+ sky130_fd_sc_hd__inv_2
Xclkbuf_2_0_0___dut__.__uuf__.__clk_source__ clkbuf_2_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1642_ __dut__.__uuf__._1642_/A VGND VGND VPWR VPWR __dut__.__uuf__._1642_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1573_ __dut__.__uuf__._1573_/A VGND VGND VPWR VPWR __dut__.__uuf__._1573_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1581__A2 mc[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2125_ __dut__.__uuf__._2138_/CLK __dut__._1239_/X __dut__.__uuf__._1342_/X
+ VGND VGND VPWR VPWR __dut__._1240_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2056_ __dut__.__uuf__._2065_/CLK __dut__._1101_/X __dut__.__uuf__._1598_/X
+ VGND VGND VPWR VPWR __dut__._1102_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1097__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1123_ __dut__._1129_/A1 __dut__._1123_/A2 __dut__._1122_/X VGND VGND VPWR
+ VPWR __dut__._1123_/X sky130_fd_sc_hd__a21o_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1054_ __dut__._1054_/A __dut__._1054_/B VGND VGND VPWR VPWR __dut__._1054_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1909_ __dut__._0869_/X VGND VGND VPWR VPWR __dut__.__uuf__._1914_/B
+ sky130_fd_sc_hd__inv_2
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1021__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0907_ __dut__._1383_/A1 prod[50] __dut__._0906_/X VGND VGND VPWR VPWR __dut__._1870_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1887_ clkbuf_4_9_0_tck/X __dut__._1887_/D __dut__._1442_/Y VGND VGND VPWR
+ VPWR __dut__._1887_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1823__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1079__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1214__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1251__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1625_ __dut__.__uuf__._1637_/A VGND VGND VPWR VPWR __dut__.__uuf__._1630_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1810_ clkbuf_4_6_0_tck/X __dut__._1810_/D __dut__._1519_/Y VGND VGND VPWR
+ VPWR __dut__._1810_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1556_ __dut__.__uuf__._1720_/A VGND VGND VPWR VPWR __dut__.__uuf__._1660_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1487_ __dut__.__uuf__._1551_/A VGND VGND VPWR VPWR __dut__.__uuf__._1487_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1741_ __dut__._1543_/Y mp[22] __dut__._1740_/X VGND VGND VPWR VPWR __dut__._1741_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1672_ __dut__._1788_/A __dut__._1822_/Q VGND VGND VPWR VPWR __dut__._1672_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1846__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2108_ __dut__.__uuf__._2208_/CLK __dut__._1205_/X __dut__.__uuf__._1428_/X
+ VGND VGND VPWR VPWR __dut__._1206_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2039_ __dut__.__uuf__._2083_/CLK __dut__._1067_/X __dut__.__uuf__._1620_/X
+ VGND VGND VPWR VPWR __dut__._1068_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_51_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1106_ __dut__._1106_/A __dut__._1106_/B VGND VGND VPWR VPWR __dut__._1106_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1037_ __dut__._1037_/A1 __dut__._1037_/A2 __dut__._1036_/X VGND VGND VPWR
+ VPWR __dut__._1037_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1545__A2 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2107__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_90_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_113_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1233__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__292__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1410_ __dut__._1216_/B VGND VGND VPWR VPWR __dut__.__uuf__._1410_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1341_ __dut__.__uuf__._1329_/X __dut__.__uuf__._1339_/X __dut__._1242_/B
+ __dut__.__uuf__._1340_/X VGND VGND VPWR VPWR __dut__._1241_/A2 sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._1869__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1272_ __dut__.__uuf__._1267_/Y __dut__.__uuf__._2004_/B __dut__.__uuf__._1271_/X
+ VGND VGND VPWR VPWR __dut__._1267_/A2 sky130_fd_sc_hd__o21ai_4
XFILLER_100_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_5 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1389_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__309__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1608_ __dut__.__uuf__._1611_/A VGND VGND VPWR VPWR __dut__.__uuf__._1608_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1539_ __dut__.__uuf__._1530_/X __dut__.__uuf__._1526_/X __dut__._1158_/B
+ __dut__.__uuf__._1535_/X __dut__.__uuf__._1538_/X VGND VGND VPWR VPWR __dut__._1157_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1724_ __dut__._1788_/A __dut__._1835_/Q VGND VGND VPWR VPWR __dut__._1724_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_99_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1655_ __dut__._1655_/A1 __dut__._1653_/X __dut__._1654_/X VGND VGND VPWR
+ VPWR __dut__._1817_/D sky130_fd_sc_hd__a21o_4
X__dut__._1586_ __dut__._1766_/A __dut__._1799_/Q VGND VGND VPWR VPWR __dut__._1586_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._0958__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1215__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0868__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1890_ __dut__.__uuf__._1890_/A VGND VGND VPWR VPWR __dut__._1089_/A2
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1757__A2 mp[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_12 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0983_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_45 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._1331_/A1
+ sky130_fd_sc_hd__buf_4
Xpsn_inst_psn_buff_56 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1735_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_34 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._0961_/A1
+ sky130_fd_sc_hd__buf_4
Xpsn_inst_psn_buff_23 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0943_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_78 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1129_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_67 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1651_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_89 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1273_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1324_ __dut__.__uuf__._1324_/A VGND VGND VPWR VPWR __dut__.__uuf__._1324_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1255_ __dut__.__uuf__._1242_/X __dut__.__uuf__._1254_/X prod[4]
+ prod[5] __dut__.__uuf__._1249_/X VGND VGND VPWR VPWR __dut__._1277_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_86_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1186_ __dut__.__uuf__._1183_/X __dut__.__uuf__._1180_/X prod[27]
+ prod[28] __dut__.__uuf__._1175_/X VGND VGND VPWR VPWR __dut__._1323_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1693__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1440_ rst VGND VGND VPWR VPWR __dut__._1440_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1371_ __dut__._1383_/A1 __dut__._1371_/A2 __dut__._1370_/X VGND VGND VPWR
+ VPWR __dut__._1371_/X sky130_fd_sc_hd__a21o_4
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1402__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_250_ _199_/X _314_/Q VGND VGND VPWR VPWR _250_/Q sky130_fd_sc_hd__dfxtp_4
X_181_ _271_/Q _182_/B VGND VGND VPWR VPWR _270_/D sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_14_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1707_ __dut__._1719_/A1 __dut__._1705_/X __dut__._1706_/X VGND VGND VPWR
+ VPWR __dut__._1830_/D sky130_fd_sc_hd__a21o_4
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1638_ __dut__._1638_/A __dut__._1811_/Q VGND VGND VPWR VPWR __dut__._1638_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1569_ __dut__._1543_/Y mc[15] __dut__._1568_/X VGND VGND VPWR VPWR __dut__._1569_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_1_0___dut__.__uuf__.__clk_source__ clkbuf_4_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2049_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1675__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1040_ __dut__.__uuf__._1190_/A __dut__.__uuf__._1295_/A VGND VGND
+ VPWR VPWR __dut__.__uuf__._1448_/A sky130_fd_sc_hd__or2_4
XFILLER_83_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1907__CLK __dut__._1919_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1942_ __dut__._1765_/X VGND VGND VPWR VPWR __dut__.__uuf__._1948_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_24_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1873_ __dut__._1086_/B VGND VGND VPWR VPWR __dut__.__uuf__._1873_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1222__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0940_ __dut__._0940_/A __dut__._1886_/Q VGND VGND VPWR VPWR __dut__._0940_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._0871_ __dut__._1767_/A1 __dut__._0869_/X __dut__._0870_/X VGND VGND VPWR
+ VPWR __dut__._1853_/D sky130_fd_sc_hd__a21o_4
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1307_ __dut__.__uuf__._1316_/A VGND VGND VPWR VPWR __dut__.__uuf__._1307_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_59_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1238_ __dut__.__uuf__._1450_/A VGND VGND VPWR VPWR __dut__.__uuf__._1483_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1423_ rst VGND VGND VPWR VPWR __dut__._1423_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1169_ __dut__.__uuf__._1168_/X __dut__.__uuf__._1165_/X prod[33]
+ prod[34] __dut__.__uuf__._1160_/X VGND VGND VPWR VPWR __dut__._1335_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1354_ __dut__._1378_/A prod[42] VGND VGND VPWR VPWR __dut__._1354_/X sky130_fd_sc_hd__and2_4
XFILLER_27_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1285_ __dut__._1285_/A1 __dut__._1285_/A2 __dut__._1284_/X VGND VGND VPWR
+ VPWR __dut__._1285_/X sky130_fd_sc_hd__a21o_4
XFILLER_30_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_302_ _194_/A _302_/D trst VGND VGND VPWR VPWR _302_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1132__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_233_ _291_/Q _298_/Q _305_/Q _306_/Q VGND VGND VPWR VPWR _234_/B sky130_fd_sc_hd__or4_4
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_164_ _285_/Q _164_/B VGND VGND VPWR VPWR _284_/D sky130_fd_sc_hd__and2_4
XFILLER_69_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1657__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2210_ __dut__.__uuf__._2210_/CLK __dut__._1409_/X __dut__.__uuf__._2008_/X
+ VGND VGND VPWR VPWR __dut__._0936_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__279__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2141_ __dut__.__uuf__._2208_/CLK __dut__._1271_/X __dut__.__uuf__._1261_/X
+ VGND VGND VPWR VPWR prod[1] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2072_ __dut__.__uuf__._2114_/CLK __dut__._1133_/X __dut__.__uuf__._1578_/X
+ VGND VGND VPWR VPWR __dut__._1134_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_96_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1023_ __dut__.__uuf__._2005_/C VGND VGND VPWR VPWR __dut__.__uuf__._1024_/C
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._0871__A2 __dut__._0869_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1925_ __dut__.__uuf__._1968_/A __dut__.__uuf__._1925_/B __dut__.__uuf__._1925_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1927_/B sky130_fd_sc_hd__or3_4
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1070_ __dut__._1074_/A __dut__._1070_/B VGND VGND VPWR VPWR __dut__._1070_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1856_ __dut__.__uuf__._1851_/Y __dut__.__uuf__._1852_/Y __dut__.__uuf__._1831_/X
+ __dut__.__uuf__._1855_/X VGND VGND VPWR VPWR __dut__.__uuf__._1857_/A sky130_fd_sc_hd__a211o_4
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1787_ __dut__._1048_/B VGND VGND VPWR VPWR __dut__.__uuf__._1787_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._0923_ __dut__._1383_/A1 prod[58] __dut__._0922_/X VGND VGND VPWR VPWR __dut__._1878_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_86_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_81_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1639__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1406_ __dut__._1408_/A __dut__._1406_/B VGND VGND VPWR VPWR __dut__._1406_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1337_ __dut__._1339_/A1 __dut__._1337_/A2 __dut__._1336_/X VGND VGND VPWR
+ VPWR __dut__._1337_/X sky130_fd_sc_hd__a21o_4
XFILLER_74_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2140__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1268_ __dut__._1786_/A __dut__._1268_/B VGND VGND VPWR VPWR __dut__._1268_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1199_ __dut__._1779_/A1 __dut__._1199_/A2 __dut__._1198_/X VGND VGND VPWR
+ VPWR __dut__._1199_/X sky130_fd_sc_hd__a21o_4
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_216_ _294_/Q _292_/Q _232_/A VGND VGND VPWR VPWR _291_/D sky130_fd_sc_hd__o21a_4
X_147_ _310_/Q _239_/A VGND VGND VPWR VPWR _147_/X sky130_fd_sc_hd__and2_4
XFILLER_93_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_143_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1710_ __dut__.__uuf__._1706_/Y __dut__.__uuf__._1707_/Y __dut__.__uuf__._1660_/X
+ __dut__.__uuf__._1709_/X VGND VGND VPWR VPWR __dut__.__uuf__._1711_/A sky130_fd_sc_hd__a211o_4
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1641_ __dut__.__uuf__._1642_/A VGND VGND VPWR VPWR __dut__.__uuf__._1641_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1500__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1572_ __dut__.__uuf__._1908_/A VGND VGND VPWR VPWR __dut__.__uuf__._1573_/A
+ sky130_fd_sc_hd__buf_2
Xclkbuf_2_0_0_tck clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR clkbuf_3_1_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2124_ __dut__.__uuf__._2138_/CLK __dut__._1237_/X __dut__.__uuf__._1347_/X
+ VGND VGND VPWR VPWR __dut__._1238_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._2013__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2055_ __dut__.__uuf__._2065_/CLK __dut__._1099_/X __dut__.__uuf__._1599_/X
+ VGND VGND VPWR VPWR __dut__._1100_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2163__CLK __dut__.__uuf__._2164_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1122_ __dut__._1678_/A __dut__._1122_/B VGND VGND VPWR VPWR __dut__._1122_/X
+ sky130_fd_sc_hd__and2_4
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1053_ __dut__._1053_/A1 __dut__._1053_/A2 __dut__._1052_/X VGND VGND VPWR
+ VPWR __dut__._1053_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1908_ __dut__.__uuf__._1908_/A VGND VGND VPWR VPWR __dut__.__uuf__._1908_/X
+ sky130_fd_sc_hd__buf_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1839_ __dut__.__uuf__._1826_/X __dut__.__uuf__._1838_/B __dut__.__uuf__._1838_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1840_/C sky130_fd_sc_hd__o21ai_4
XANTENNA___dut__._1410__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0906_ __dut__._1378_/A __dut__._1869_/Q VGND VGND VPWR VPWR __dut__._0906_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_4_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1886_ clkbuf_4_9_0_tck/X __dut__._1886_/D __dut__._1443_/Y VGND VGND VPWR
+ VPWR __dut__._1886_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1320__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2036__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1887__A __dut__._1549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1798__CLK __dut__._1410_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1230__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1624_ __dut__.__uuf__._1624_/A VGND VGND VPWR VPWR __dut__.__uuf__._1624_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1555_ __dut__.__uuf__._1569_/A VGND VGND VPWR VPWR __dut__.__uuf__._1555_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1740_ __dut__._1788_/A __dut__._1839_/Q VGND VGND VPWR VPWR __dut__._1740_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1486_ __dut__.__uuf__._1486_/A VGND VGND VPWR VPWR __dut__.__uuf__._1486_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1671_ __dut__._1767_/A1 __dut__._1669_/X __dut__._1670_/X VGND VGND VPWR
+ VPWR __dut__._1821_/D sky130_fd_sc_hd__a21o_4
XFILLER_88_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2107_ __dut__.__uuf__._2107_/CLK __dut__._1203_/X __dut__.__uuf__._1432_/X
+ VGND VGND VPWR VPWR __dut__._1204_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_67_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2038_ __dut__.__uuf__._2083_/CLK __dut__._1065_/X __dut__.__uuf__._1621_/X
+ VGND VGND VPWR VPWR __dut__._1066_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_44_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1105_ __dut__._1129_/A1 __dut__._1105_/A2 __dut__._1104_/X VGND VGND VPWR
+ VPWR __dut__._1105_/X sky130_fd_sc_hd__a21o_4
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1036_ __dut__._1678_/A __dut__._1036_/B VGND VGND VPWR VPWR __dut__._1036_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1869_ __dut__._1915_/CLK __dut__._1869_/D __dut__._1460_/Y VGND VGND VPWR
+ VPWR __dut__._1869_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_95_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_106_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1050__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1340_ __dut__.__uuf__._1380_/A VGND VGND VPWR VPWR __dut__.__uuf__._1340_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1271_ __dut__.__uuf__._1401_/A VGND VGND VPWR VPWR __dut__.__uuf__._1271_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_85_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2201__CLK __dut__.__uuf__._2210_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_6 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0883_/A1 sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1607_ __dut__.__uuf__._1611_/A VGND VGND VPWR VPWR __dut__.__uuf__._1607_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1538_ __dut__._1681_/X __dut__.__uuf__._1536_/X __dut__._1160_/B
+ __dut__.__uuf__._1537_/X VGND VGND VPWR VPWR __dut__.__uuf__._1538_/X sky130_fd_sc_hd__o22a_4
X__dut__._1723_ __dut__._1767_/A1 __dut__._1721_/X __dut__._1722_/X VGND VGND VPWR
+ VPWR __dut__._1834_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1469_ __dut__.__uuf__._1469_/A VGND VGND VPWR VPWR __dut__.__uuf__._1486_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1654_ __dut__._1766_/A __dut__._1816_/Q VGND VGND VPWR VPWR __dut__._1654_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1585_ __dut__._1543_/Y mc[19] __dut__._1584_/X VGND VGND VPWR VPWR __dut__._1585_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1019_ __dut__._1129_/A1 __dut__._1019_/A2 __dut__._1018_/X VGND VGND VPWR
+ VPWR __dut__._1019_/X sky130_fd_sc_hd__a21o_4
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0884__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_13 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0981_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1836__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_46 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._1323_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_35 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._1291_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_24 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1277_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_68 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1679_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_79 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1647_/A1
+ sky130_fd_sc_hd__buf_4
Xpsn_inst_psn_buff_57 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1731_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1323_ __dut__.__uuf__._1400_/A VGND VGND VPWR VPWR __dut__.__uuf__._1323_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1254_ __dut__.__uuf__._1483_/A VGND VGND VPWR VPWR __dut__.__uuf__._1254_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1185_ __dut__.__uuf__._1189_/A VGND VGND VPWR VPWR __dut__.__uuf__._1185_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1693__A2 mp[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1370_ __dut__._1378_/A prod[50] VGND VGND VPWR VPWR __dut__._1370_/X sky130_fd_sc_hd__and2_4
XFILLER_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_180_ _272_/Q _187_/B VGND VGND VPWR VPWR _271_/D sky130_fd_sc_hd__or2_4
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1381__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1706_ __dut__._1766_/A __dut__._1829_/Q VGND VGND VPWR VPWR __dut__._1706_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1133__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1637_ __dut__._1543_/Y mc[30] __dut__._1636_/X VGND VGND VPWR VPWR __dut__._1637_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1568_ __dut__._1788_/A __dut__._1796_/Q VGND VGND VPWR VPWR __dut__._1568_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1499_ rst VGND VGND VPWR VPWR __dut__._1499_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_173_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1941_ __dut__.__uuf__._1941_/A VGND VGND VPWR VPWR __dut__.__uuf__._1941_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1872_ __dut__.__uuf__._1883_/A __dut__.__uuf__._1872_/B __dut__.__uuf__._1872_/C
+ VGND VGND VPWR VPWR __dut__._1079_/A2 sky130_fd_sc_hd__and3_4
XANTENNA___dut__._1503__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1262__A3 prod[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0870_ __dut__._1766_/A __dut__._1852_/Q VGND VGND VPWR VPWR __dut__._0870_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1363__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2210_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1306_ __dut__.__uuf__._1303_/X __dut__.__uuf__._1305_/X __dut__._1256_/B
+ __dut__.__uuf__._1303_/X VGND VGND VPWR VPWR __dut__._1255_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1115__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1237_ __dut__.__uuf__._1248_/A VGND VGND VPWR VPWR __dut__.__uuf__._1237_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1168_ __dut__.__uuf__._1212_/A VGND VGND VPWR VPWR __dut__.__uuf__._1168_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1422_ rst VGND VGND VPWR VPWR __dut__._1422_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1099_ __dut__.__uuf__._1099_/A VGND VGND VPWR VPWR __dut__.__uuf__._1099_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1353_ __dut__._1383_/A1 __dut__._1353_/A2 __dut__._1352_/X VGND VGND VPWR
+ VPWR __dut__._1353_/X sky130_fd_sc_hd__a21o_4
X__dut__._1284_ __dut__._1770_/A prod[7] VGND VGND VPWR VPWR __dut__._1284_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1413__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_301_ _194_/A _301_/D trst VGND VGND VPWR VPWR _301_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1045__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1132__B __dut__._1132_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_232_ _232_/A _232_/B VGND VGND VPWR VPWR _304_/D sky130_fd_sc_hd__and2_4
X_163_ _286_/Q _172_/B VGND VGND VPWR VPWR _285_/D sky130_fd_sc_hd__or2_4
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0999_ __dut__._1331_/A1 prod[31] __dut__._0998_/X VGND VGND VPWR VPWR __dut__._1916_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_97_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1657__A2 mp[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1593__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2140_ __dut__.__uuf__._2208_/CLK __dut__._1269_/X __dut__.__uuf__._1263_/X
+ VGND VGND VPWR VPWR prod[0] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2071_ __dut__.__uuf__._2107_/CLK __dut__._1131_/X __dut__.__uuf__._1579_/X
+ VGND VGND VPWR VPWR __dut__._1132_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1022_ __dut__._1402_/B __dut__.__uuf__._1029_/A __dut__._1398_/B
+ __dut__.__uuf__._1022_/D VGND VGND VPWR VPWR __dut__.__uuf__._2005_/C sky130_fd_sc_hd__or4_4
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1924_ __dut__.__uuf__._1917_/Y __dut__.__uuf__._1918_/Y __dut__.__uuf__._1917_/Y
+ __dut__.__uuf__._1918_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1925_/C sky130_fd_sc_hd__a2bb2o_4
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1855_ __dut__.__uuf__._1851_/Y __dut__.__uuf__._1852_/Y __dut__.__uuf__._1853_/X
+ __dut__.__uuf__._1859_/B VGND VGND VPWR VPWR __dut__.__uuf__._1855_/X sky130_fd_sc_hd__o22a_4
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1786_ __dut__._1054_/B VGND VGND VPWR VPWR __dut__.__uuf__._1786_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_20_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._0922_ __dut__._1542_/A __dut__._1877_/Q VGND VGND VPWR VPWR __dut__._0922_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2092__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1405_ __dut__._1405_/A1 __dut__._1405_/A2 __dut__._1404_/X VGND VGND VPWR
+ VPWR __dut__._1405_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_74_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1336_ __dut__._1378_/A prod[33] VGND VGND VPWR VPWR __dut__._1336_/X sky130_fd_sc_hd__and2_4
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1267_ __dut__._1787_/A1 __dut__._1267_/A2 __dut__._1266_/X VGND VGND VPWR
+ VPWR __dut__._1267_/X sky130_fd_sc_hd__a21o_4
X__dut__._1198_ __dut__._1198_/A __dut__._1198_/B VGND VGND VPWR VPWR __dut__._1198_/X
+ sky130_fd_sc_hd__and2_4
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1575__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_215_ _225_/B VGND VGND VPWR VPWR _232_/A sky130_fd_sc_hd__buf_2
XFILLER_7_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_146_ _239_/A VGND VGND VPWR VPWR _146_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_136_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._0892__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1640_ __dut__.__uuf__._1642_/A VGND VGND VPWR VPWR __dut__.__uuf__._1640_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1571_ __dut__.__uuf__._1685_/A VGND VGND VPWR VPWR __dut__.__uuf__._1908_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_88_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1228__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2123_ __dut__.__uuf__._2138_/CLK __dut__._1235_/X __dut__.__uuf__._1353_/X
+ VGND VGND VPWR VPWR __dut__._1236_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2054_ __dut__.__uuf__._2065_/CLK __dut__._1097_/X __dut__.__uuf__._1601_/X
+ VGND VGND VPWR VPWR __dut__._1098_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_29_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1121_ __dut__._1129_/A1 __dut__._1121_/A2 __dut__._1120_/X VGND VGND VPWR
+ VPWR __dut__._1121_/X sky130_fd_sc_hd__a21o_4
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1052_ __dut__._1678_/A __dut__._1052_/B VGND VGND VPWR VPWR __dut__._1052_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1907_ __dut__._1092_/B VGND VGND VPWR VPWR __dut__.__uuf__._1907_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1838_ __dut__.__uuf__._1859_/A __dut__.__uuf__._1838_/B __dut__.__uuf__._1838_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1840_/B sky130_fd_sc_hd__or3_4
XANTENNA___dut__._1557__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1410__B __dut__._1410_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1769_ __dut__.__uuf__._1763_/Y __dut__.__uuf__._1764_/Y __dut__.__uuf__._1763_/Y
+ __dut__.__uuf__._1764_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1770_/C sky130_fd_sc_hd__a2bb2o_4
X__dut__._0905_ __dut__._1383_/A1 prod[49] __dut__._0904_/X VGND VGND VPWR VPWR __dut__._1869_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1885_ clkbuf_4_9_0_tck/X __dut__._1885_/D __dut__._1444_/Y VGND VGND VPWR
+ VPWR __dut__._1885_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_psn_inst_psn_buff_8_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1319_ __dut__._1319_/A1 __dut__._1319_/A2 __dut__._1318_/X VGND VGND VPWR
+ VPWR __dut__._1319_/X sky130_fd_sc_hd__a21o_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__269__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_129_ _121_/Y _231_/A _125_/X _128_/X VGND VGND VPWR VPWR _130_/A sky130_fd_sc_hd__a211o_4
XFILLER_98_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1048__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1787__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1511__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1623_ __dut__.__uuf__._1624_/A VGND VGND VPWR VPWR __dut__.__uuf__._1623_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1554_ __dut__.__uuf__._1575_/A VGND VGND VPWR VPWR __dut__.__uuf__._1569_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1485_ __dut__.__uuf__._1466_/X __dut__.__uuf__._1483_/X __dut__._1182_/B
+ __dut__.__uuf__._1471_/X __dut__.__uuf__._1484_/X VGND VGND VPWR VPWR __dut__._1181_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1670_ __dut__._1766_/A __dut__._1820_/Q VGND VGND VPWR VPWR __dut__._1670_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2106_ __dut__.__uuf__._2208_/CLK __dut__._1201_/X __dut__.__uuf__._1436_/X
+ VGND VGND VPWR VPWR __dut__._1202_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2037_ __dut__.__uuf__._2083_/CLK __dut__._1063_/X __dut__.__uuf__._1622_/X
+ VGND VGND VPWR VPWR __dut__._1064_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1104_ __dut__._1678_/A __dut__._1104_/B VGND VGND VPWR VPWR __dut__._1104_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1421__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1035_ __dut__._1129_/A1 __dut__._1035_/A2 __dut__._1034_/X VGND VGND VPWR
+ VPWR __dut__._1035_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_37_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1892__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1868_ __dut__._1915_/CLK __dut__._1868_/D __dut__._1461_/Y VGND VGND VPWR
+ VPWR __dut__._1868_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1799_ __dut__._1410_/B __dut__._1799_/D __dut__._1530_/Y VGND VGND VPWR
+ VPWR __dut__._1799_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1769__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._1898__A __dut__._0873_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1270_ __dut__._1781_/X __dut__.__uuf__._1295_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1401_/A sky130_fd_sc_hd__nand2_4
XFILLER_98_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1506__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_7 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0881_/A1 sky130_fd_sc_hd__buf_2
XFILLER_22_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1044__A1 __dut__.__uuf__._1100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1606_ __dut__.__uuf__._1606_/A VGND VGND VPWR VPWR __dut__.__uuf__._1611_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1537_ __dut__.__uuf__._1720_/A VGND VGND VPWR VPWR __dut__.__uuf__._1537_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_1_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1722_ __dut__._1766_/A __dut__._1823_/Q VGND VGND VPWR VPWR __dut__._1722_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1468_ __dut__.__uuf__._1466_/X __dut__.__uuf__._1462_/X __dut__._1190_/B
+ __dut__.__uuf__._1449_/X __dut__.__uuf__._1467_/X VGND VGND VPWR VPWR __dut__._1189_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1653_ __dut__._1543_/Y mp[2] __dut__._1652_/X VGND VGND VPWR VPWR __dut__._1653_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1399_ __dut__._1220_/B VGND VGND VPWR VPWR __dut__.__uuf__._1399_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1416__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1584_ __dut__._1788_/A __dut__._1800_/Q VGND VGND VPWR VPWR __dut__._1584_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._1048__A __dut__.__uuf__._2008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1018_ __dut__._1128_/A __dut__._1018_/B VGND VGND VPWR VPWR __dut__._1018_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA__307__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1326__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_47 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._0989_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_14 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1313_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_25 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1279_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_36 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._1293_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_69 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1047_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_58 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1727_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1322_ __dut__._1250_/B VGND VGND VPWR VPWR __dut__.__uuf__._1322_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1253_ __dut__.__uuf__._1263_/A VGND VGND VPWR VPWR __dut__.__uuf__._1253_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1184_ __dut__.__uuf__._1183_/X __dut__.__uuf__._1180_/X prod[28]
+ prod[29] __dut__.__uuf__._1175_/X VGND VGND VPWR VPWR __dut__._1325_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_86_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1236__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2049__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1705_ __dut__._1543_/Y mp[14] __dut__._1704_/X VGND VGND VPWR VPWR __dut__._1705_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1636_ __dut__._1788_/A __dut__._1813_/Q VGND VGND VPWR VPWR __dut__._1636_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1567_ __dut__._1767_/A1 __dut__._1565_/X __dut__._1566_/X VGND VGND VPWR
+ VPWR __dut__._1795_/D sky130_fd_sc_hd__a21o_4
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1498_ rst VGND VGND VPWR VPWR __dut__._1498_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_166_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1803__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1940_ __dut__._1104_/B VGND VGND VPWR VPWR __dut__.__uuf__._1940_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1871_ __dut__.__uuf__._1826_/X __dut__.__uuf__._1870_/B __dut__.__uuf__._1870_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1872_/C sky130_fd_sc_hd__o21ai_4
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1305_ __dut__.__uuf__._1304_/Y __dut__.__uuf__._1297_/X __dut__.__uuf__._1299_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1305_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_3_3_0___dut__.__uuf__.__clk_source__ clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_7_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1236_ __dut__.__uuf__._1236_/A VGND VGND VPWR VPWR __dut__.__uuf__._1248_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1167_ __dut__.__uuf__._1174_/A VGND VGND VPWR VPWR __dut__.__uuf__._1167_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1421_ rst VGND VGND VPWR VPWR __dut__._1421_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1098_ __dut__.__uuf__._1093_/X __dut__.__uuf__._1090_/X prod[56]
+ prod[57] __dut__.__uuf__._1085_/X VGND VGND VPWR VPWR __dut__._1381_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1352_ __dut__._1378_/A prod[41] VGND VGND VPWR VPWR __dut__._1352_/X sky130_fd_sc_hd__and2_4
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1283_ __dut__._1283_/A1 __dut__._1283_/A2 __dut__._1282_/X VGND VGND VPWR
+ VPWR __dut__._1283_/X sky130_fd_sc_hd__a21o_4
X_300_ _194_/A _300_/D trst VGND VGND VPWR VPWR _300_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_91_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._0929__A2 prod[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_231_ _231_/A _298_/Q _305_/Q VGND VGND VPWR VPWR _232_/B sky130_fd_sc_hd__or3_4
XANTENNA___dut__._1051__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_162_ _287_/Q _164_/B VGND VGND VPWR VPWR _286_/D sky130_fd_sc_hd__and2_4
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._0998_ __dut__._1378_/A __dut__._1915_/Q VGND VGND VPWR VPWR __dut__._0998_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1619_ __dut__._1767_/A1 __dut__._1617_/X __dut__._1618_/X VGND VGND VPWR
+ VPWR __dut__._1808_/D sky130_fd_sc_hd__a21o_4
XFILLER_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0865__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1604__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1593__A2 mc[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2070_ __dut__.__uuf__._2107_/CLK __dut__._1129_/X __dut__.__uuf__._1580_/X
+ VGND VGND VPWR VPWR __dut__._1130_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1021_ __dut__.__uuf__._1036_/A __dut__._1408_/B __dut__._1406_/B
+ __dut__._1404_/B VGND VGND VPWR VPWR __dut__.__uuf__._1022_/D sky130_fd_sc_hd__or4_4
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1514__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1923_ __dut__.__uuf__._1923_/A VGND VGND VPWR VPWR __dut__.__uuf__._1968_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1854_ __dut__._1561_/X VGND VGND VPWR VPWR __dut__.__uuf__._1859_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1033__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1785_ __dut__.__uuf__._1828_/A __dut__.__uuf__._1785_/B __dut__.__uuf__._1785_/C
+ VGND VGND VPWR VPWR __dut__._1047_/A2 sky130_fd_sc_hd__and3_4
X__dut__._0921_ __dut__._0921_/A1 prod[57] __dut__._0920_/X VGND VGND VPWR VPWR __dut__._1877_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1849__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1219_ __dut__.__uuf__._1249_/A VGND VGND VPWR VPWR __dut__.__uuf__._1219_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2199_ __dut__.__uuf__._2200_/CLK __dut__._1387_/X __dut__.__uuf__._1088_/X
+ VGND VGND VPWR VPWR prod[59] sky130_fd_sc_hd__dfrtp_4
XFILLER_74_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1404_ __dut__._1404_/A __dut__._1404_/B VGND VGND VPWR VPWR __dut__._1404_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1335_ __dut__._1339_/A1 __dut__._1335_/A2 __dut__._1334_/X VGND VGND VPWR
+ VPWR __dut__._1335_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1424__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_67_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1266_ __dut__._1786_/A __dut__._1266_/B VGND VGND VPWR VPWR __dut__._1266_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1197_ __dut__._1197_/A1 __dut__._1197_/A2 __dut__._1196_/X VGND VGND VPWR
+ VPWR __dut__._1197_/X sky130_fd_sc_hd__a21o_4
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ _234_/A _214_/B VGND VGND VPWR VPWR _225_/B sky130_fd_sc_hd__nor2_4
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_145_ _239_/A _142_/Y tdi _310_/Q _144_/Y VGND VGND VPWR VPWR _310_/D sky130_fd_sc_hd__a32o_4
XFILLER_38_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1334__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_129_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1263__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1015__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1570_ __dut__._1140_/B VGND VGND VPWR VPWR __dut__.__uuf__._1685_/A
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1509__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2122_ __dut__.__uuf__._2138_/CLK __dut__._1233_/X __dut__.__uuf__._1358_/X
+ VGND VGND VPWR VPWR __dut__._1234_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2053_ __dut__.__uuf__._2065_/CLK __dut__._1095_/X __dut__.__uuf__._1602_/X
+ VGND VGND VPWR VPWR __dut__._1096_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1244__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1120_ __dut__._1678_/A __dut__._1120_/B VGND VGND VPWR VPWR __dut__._1120_/X
+ sky130_fd_sc_hd__and2_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1051_ __dut__._1767_/A1 __dut__._1051_/A2 __dut__._1050_/X VGND VGND VPWR
+ VPWR __dut__._1051_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1906_ __dut__._1098_/B VGND VGND VPWR VPWR __dut__.__uuf__._1906_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1837_ __dut__.__uuf__._1829_/Y __dut__.__uuf__._1830_/Y __dut__.__uuf__._1829_/Y
+ __dut__.__uuf__._1830_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1838_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._1557__A2 mc[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1768_ __dut__.__uuf__._1768_/A VGND VGND VPWR VPWR __dut__._1045_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1699_ __dut__.__uuf__._1695_/Y __dut__.__uuf__._1696_/Y __dut__.__uuf__._1660_/X
+ __dut__.__uuf__._1698_/X VGND VGND VPWR VPWR __dut__.__uuf__._1700_/A sky130_fd_sc_hd__a211o_4
X__dut__._0904_ __dut__._1378_/A __dut__._1868_/Q VGND VGND VPWR VPWR __dut__._0904_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1884_ _290_/CLK __dut__._1884_/D __dut__._1445_/Y VGND VGND VPWR VPWR _210_/A2
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1419__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1154__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1245__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1318_ __dut__._1318_/A prod[24] VGND VGND VPWR VPWR __dut__._1318_/X sky130_fd_sc_hd__and2_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1249_ __dut__._1787_/A1 __dut__._1249_/A2 __dut__._1248_/X VGND VGND VPWR
+ VPWR __dut__._1249_/X sky130_fd_sc_hd__a21o_4
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_128_ _214_/B VGND VGND VPWR VPWR _128_/X sky130_fd_sc_hd__buf_2
XFILLER_97_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1622_ __dut__.__uuf__._1624_/A VGND VGND VPWR VPWR __dut__.__uuf__._1622_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1071__A2 __dut__.__uuf__._1069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1553_ __dut__.__uuf__._1551_/X __dut__.__uuf__._1547_/X __dut__._1150_/B
+ __dut__.__uuf__._1535_/X __dut__.__uuf__._1552_/X VGND VGND VPWR VPWR __dut__._1149_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1484_ __dut__._1733_/X __dut__.__uuf__._1472_/X __dut__._1184_/B
+ __dut__.__uuf__._1473_/X VGND VGND VPWR VPWR __dut__.__uuf__._1484_/X sky130_fd_sc_hd__o22a_4
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2105_ __dut__.__uuf__._2208_/CLK __dut__._1199_/X __dut__.__uuf__._1442_/X
+ VGND VGND VPWR VPWR __dut__._1200_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_96_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2036_ __dut__.__uuf__._2083_/CLK __dut__._1061_/X __dut__.__uuf__._1623_/X
+ VGND VGND VPWR VPWR __dut__._1062_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1227__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1103_ __dut__._1129_/A1 __dut__._1103_/A2 __dut__._1102_/X VGND VGND VPWR
+ VPWR __dut__._1103_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1702__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1034_ __dut__._1078_/A __dut__._1034_/B VGND VGND VPWR VPWR __dut__._1034_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1867_ __dut__._1915_/CLK __dut__._1867_/D __dut__._1462_/Y VGND VGND VPWR
+ VPWR __dut__._1867_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0988__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1798_ __dut__._1410_/B __dut__._1798_/D __dut__._1531_/Y VGND VGND VPWR
+ VPWR __dut__._1798_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1509__A __dut__.__uuf__._1551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1612__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1769__A2 mp[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0898__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1209__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1522__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_8 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1343_/A1 sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1605_ __dut__.__uuf__._1605_/A VGND VGND VPWR VPWR __dut__.__uuf__._1605_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1536_ __dut__.__uuf__._1536_/A VGND VGND VPWR VPWR __dut__.__uuf__._1536_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1721_ __dut__._1543_/Y mc[4] __dut__._1720_/X VGND VGND VPWR VPWR __dut__._1721_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1467_ __dut__._1749_/X __dut__.__uuf__._1451_/X __dut__._1192_/B
+ __dut__.__uuf__._1452_/X VGND VGND VPWR VPWR __dut__.__uuf__._1467_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1652_ __dut__._1788_/A __dut__._1817_/Q VGND VGND VPWR VPWR __dut__._1652_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA__259__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1398_ __dut__.__uuf__._1418_/A VGND VGND VPWR VPWR __dut__.__uuf__._1398_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_76_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1583_ __dut__._1767_/A1 __dut__._1581_/X __dut__._1582_/X VGND VGND VPWR
+ VPWR __dut__._1799_/D sky130_fd_sc_hd__a21o_4
XFILLER_72_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2019_ __dut__.__uuf__._2049_/CLK __dut__._1027_/X __dut__.__uuf__._1644_/X
+ VGND VGND VPWR VPWR __dut__._1028_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1432__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1017_ __dut__._1129_/A1 __dut__._1017_/A2 __dut__._1016_/X VGND VGND VPWR
+ VPWR __dut__._1017_/X sky130_fd_sc_hd__a21o_4
XFILLER_40_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1919_ __dut__._1919_/CLK __dut__._1919_/D __dut__._1540_/Y VGND VGND VPWR
+ VPWR __dut__._1919_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1611__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_111_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_170 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1150_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_15 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0979_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_26 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1281_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_37 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._1295_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_48 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._1319_/A1
+ sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_59 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1167_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1321_ __dut__.__uuf__._1342_/A VGND VGND VPWR VPWR __dut__.__uuf__._1321_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1252_ __dut__.__uuf__._1346_/A VGND VGND VPWR VPWR __dut__.__uuf__._1263_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_98_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1517__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1183_ __dut__.__uuf__._1212_/A VGND VGND VPWR VPWR __dut__.__uuf__._1183_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_82_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1612__A __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1519_ __dut__.__uuf__._1529_/A VGND VGND VPWR VPWR __dut__.__uuf__._1519_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1704_ __dut__._1788_/A __dut__._1830_/Q VGND VGND VPWR VPWR __dut__._1704_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1669__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1427__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_97_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1635_ __dut__._1647_/A1 __dut__._1633_/X __dut__._1634_/X VGND VGND VPWR
+ VPWR __dut__._1812_/D sky130_fd_sc_hd__a21o_4
X__dut__._1566_ __dut__._1766_/A __dut__._1794_/Q VGND VGND VPWR VPWR __dut__._1566_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_18_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1497_ rst VGND VGND VPWR VPWR __dut__._1497_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1162__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2143__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_159_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1870_ __dut__.__uuf__._1914_/A __dut__.__uuf__._1870_/B __dut__.__uuf__._1870_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1872_/B sky130_fd_sc_hd__or3_4
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1304_ __dut__._1258_/B VGND VGND VPWR VPWR __dut__.__uuf__._1304_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2016__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_101_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1235_ __dut__.__uuf__._1227_/X __dut__.__uuf__._1223_/X prod[10]
+ prod[11] __dut__.__uuf__._1234_/X VGND VGND VPWR VPWR __dut__._1289_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_101_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1166_ __dut__.__uuf__._1153_/X __dut__.__uuf__._1165_/X prod[34]
+ prod[35] __dut__.__uuf__._1160_/X VGND VGND VPWR VPWR __dut__._1337_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1420_ rst VGND VGND VPWR VPWR __dut__._1420_/Y sky130_fd_sc_hd__inv_2
X__dut__._1351_ __dut__._1383_/A1 __dut__._1351_/A2 __dut__._1350_/X VGND VGND VPWR
+ VPWR __dut__._1351_/X sky130_fd_sc_hd__a21o_4
XFILLER_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1097_ __dut__.__uuf__._1099_/A VGND VGND VPWR VPWR __dut__.__uuf__._1097_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_39_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1282_ __dut__._1770_/A prod[6] VGND VGND VPWR VPWR __dut__._1282_/X sky130_fd_sc_hd__and2_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_230_ _234_/A _304_/Q VGND VGND VPWR VPWR _303_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1710__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1999_ __dut__.__uuf__._1999_/A VGND VGND VPWR VPWR __dut__._1133_/A2
+ sky130_fd_sc_hd__inv_2
X_161_ _288_/Q _172_/B VGND VGND VPWR VPWR _287_/D sky130_fd_sc_hd__or2_4
XANTENNA_psn_inst_psn_buff_12_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0997_ __dut__._1331_/A1 prod[30] __dut__._0996_/X VGND VGND VPWR VPWR __dut__._1915_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0996__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1618_ __dut__._1766_/A __dut__._1807_/Q VGND VGND VPWR VPWR __dut__._1618_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA__302__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._0865__A2 mc[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1549_ __dut__._1543_/Y mc[10] __dut__._1548_/X VGND VGND VPWR VPWR __dut__._1549_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_14_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1620__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2039__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1020_ __dut__._0936_/B VGND VGND VPWR VPWR __dut__.__uuf__._1036_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1922_ __dut__.__uuf__._1922_/A VGND VGND VPWR VPWR __dut__._1101_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1853_ __dut__.__uuf__._1923_/A VGND VGND VPWR VPWR __dut__.__uuf__._1853_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1530__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1784_ __dut__.__uuf__._1771_/X __dut__.__uuf__._1783_/B __dut__.__uuf__._1783_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1785_/C sky130_fd_sc_hd__o21ai_4
X__dut__._0920_ __dut__._1542_/A __dut__._1876_/Q VGND VGND VPWR VPWR __dut__._0920_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_20_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1218_ __dut__.__uuf__._1218_/A VGND VGND VPWR VPWR __dut__.__uuf__._1218_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2198_ __dut__.__uuf__._2200_/CLK __dut__._1385_/X __dut__.__uuf__._1092_/X
+ VGND VGND VPWR VPWR prod[58] sky130_fd_sc_hd__dfrtp_4
X__dut__._1403_ __dut__._1405_/A1 __dut__._1403_/A2 __dut__._1402_/X VGND VGND VPWR
+ VPWR __dut__._1403_/X sky130_fd_sc_hd__a21o_4
XFILLER_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1149_ __dut__.__uuf__._1149_/A VGND VGND VPWR VPWR __dut__.__uuf__._1149_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1334_ __dut__._1378_/A prod[32] VGND VGND VPWR VPWR __dut__._1334_/X sky130_fd_sc_hd__and2_4
X__dut__._1265_ __dut__._1787_/A1 __dut__._1265_/A2 __dut__._1264_/X VGND VGND VPWR
+ VPWR __dut__._1265_/X sky130_fd_sc_hd__a21o_4
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1440__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1196_ __dut__._1274_/A __dut__._1196_/B VGND VGND VPWR VPWR __dut__._1196_/X
+ sky130_fd_sc_hd__and2_4
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ tms VGND VGND VPWR VPWR _234_/A sky130_fd_sc_hd__inv_2
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_144_ _220_/A VGND VGND VPWR VPWR _144_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1350__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__.__uuf__._1083__B1 prod[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__295__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2121_ __dut__.__uuf__._2138_/CLK __dut__._1231_/X __dut__.__uuf__._1362_/X
+ VGND VGND VPWR VPWR __dut__._1232_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2052_ __dut__.__uuf__._2065_/CLK __dut__._1093_/X __dut__.__uuf__._1603_/X
+ VGND VGND VPWR VPWR __dut__._1094_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1525__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2204__CLK __dut__.__uuf__._2210_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1905_ __dut__.__uuf__._1938_/A __dut__.__uuf__._1905_/B __dut__.__uuf__._1905_/C
+ VGND VGND VPWR VPWR __dut__._1091_/A2 sky130_fd_sc_hd__and3_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1050_ __dut__._1766_/A __dut__._1050_/B VGND VGND VPWR VPWR __dut__._1050_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1260__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1836_ __dut__.__uuf__._1946_/A VGND VGND VPWR VPWR __dut__.__uuf__._1883_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1767_ __dut__.__uuf__._1763_/Y __dut__.__uuf__._1764_/Y __dut__.__uuf__._1721_/X
+ __dut__.__uuf__._1766_/X VGND VGND VPWR VPWR __dut__.__uuf__._1768_/A sky130_fd_sc_hd__a211o_4
X__dut__.__uuf__._1698_ __dut__.__uuf__._1695_/Y __dut__.__uuf__._1696_/Y __dut__.__uuf__._1686_/X
+ __dut__.__uuf__._1703_/B VGND VGND VPWR VPWR __dut__.__uuf__._1698_/X sky130_fd_sc_hd__o22a_4
X__dut__._0903_ __dut__._1383_/A1 prod[48] __dut__._0902_/X VGND VGND VPWR VPWR __dut__._1868_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1883_ __dut__._1883_/CLK __dut__._1883_/D __dut__._1446_/Y VGND VGND VPWR
+ VPWR __dut__._1883_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1435__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1067__A __dut__.__uuf__._2008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1317_ __dut__._1339_/A1 __dut__._1317_/A2 __dut__._1316_/X VGND VGND VPWR
+ VPWR __dut__._1317_/X sky130_fd_sc_hd__a21o_4
XFILLER_28_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1248_ __dut__._1408_/A __dut__._1248_/B VGND VGND VPWR VPWR __dut__._1248_/X
+ sky130_fd_sc_hd__and2_4
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1179_ __dut__._1193_/A1 __dut__._1179_/A2 __dut__._1178_/X VGND VGND VPWR
+ VPWR __dut__._1179_/X sky130_fd_sc_hd__a21o_4
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_127_ tms _257_/D _258_/Q _127_/D VGND VGND VPWR VPWR _214_/B sky130_fd_sc_hd__and4_4
XANTENNA___dut__.__uuf__._1530__A __dut__.__uuf__._1551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_141_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1080__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1621_ __dut__.__uuf__._1624_/A VGND VGND VPWR VPWR __dut__.__uuf__._1621_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1839__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1552_ __dut__._1661_/X __dut__.__uuf__._1536_/X __dut__._1152_/B
+ __dut__.__uuf__._1537_/X VGND VGND VPWR VPWR __dut__.__uuf__._1552_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1483_ __dut__.__uuf__._1483_/A VGND VGND VPWR VPWR __dut__.__uuf__._1483_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2104_ __dut__.__uuf__._2208_/CLK __dut__._1197_/X __dut__.__uuf__._1447_/X
+ VGND VGND VPWR VPWR __dut__._1198_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_69_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2035_ __dut__.__uuf__._2083_/CLK __dut__._1059_/X __dut__.__uuf__._1624_/X
+ VGND VGND VPWR VPWR __dut__._1060_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1102_ __dut__._1102_/A __dut__._1102_/B VGND VGND VPWR VPWR __dut__._1102_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1033_ __dut__._1129_/A1 __dut__._1033_/A2 __dut__._1032_/X VGND VGND VPWR
+ VPWR __dut__._1033_/X sky130_fd_sc_hd__a21o_4
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1819_ __dut__._1060_/B VGND VGND VPWR VPWR __dut__.__uuf__._1819_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1866_ __dut__._1915_/CLK __dut__._1866_/D __dut__._1463_/Y VGND VGND VPWR
+ VPWR __dut__._1866_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1797_ clkbuf_4_5_0_tck/X __dut__._1797_/D __dut__._1532_/Y VGND VGND VPWR
+ VPWR __dut__._1797_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._0901__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_1_0_tck_A clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_9 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0877_/A1 sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1604_ __dut__.__uuf__._1605_/A VGND VGND VPWR VPWR __dut__.__uuf__._1604_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1535_ __dut__.__uuf__._1535_/A VGND VGND VPWR VPWR __dut__.__uuf__._1535_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1720_ __dut__._1788_/A __dut__._1834_/Q VGND VGND VPWR VPWR __dut__._1720_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1145__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1466_ __dut__.__uuf__._1466_/A VGND VGND VPWR VPWR __dut__.__uuf__._1466_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1651_ __dut__._1651_/A1 __dut__._1649_/X __dut__._1650_/X VGND VGND VPWR
+ VPWR __dut__._1816_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1397_ __dut__.__uuf__._1469_/A VGND VGND VPWR VPWR __dut__.__uuf__._1418_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1582_ __dut__._1766_/A __dut__._1798_/Q VGND VGND VPWR VPWR __dut__._1582_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2018_ __dut__.__uuf__._2049_/CLK __dut__._1025_/X __dut__.__uuf__._1645_/X
+ VGND VGND VPWR VPWR __dut__._1026_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_72_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_42_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1016_ __dut__._1128_/A __dut__._1016_/B VGND VGND VPWR VPWR __dut__._1016_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1918_ __dut__._1919_/CLK __dut__._1918_/D __dut__._1541_/Y VGND VGND VPWR
+ VPWR __dut__._1918_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2072__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1849_ _194_/A __dut__._1849_/D __dut__._1480_/Y VGND VGND VPWR VPWR __dut__._1849_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1611__A2 __dut__._1609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_160 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._0880_/A sky130_fd_sc_hd__buf_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_104_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_171 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1766_/A sky130_fd_sc_hd__buf_8
XANTENNA___dut__._1375__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_16 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1311_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_27 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0945_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_38 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._1299_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_49 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._1339_/A1
+ sky130_fd_sc_hd__buf_8
X__dut__.__uuf__._1320_ __dut__.__uuf__._1346_/A VGND VGND VPWR VPWR __dut__.__uuf__._1342_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1127__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1251_ __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR __dut__.__uuf__._1346_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1182_ __dut__.__uuf__._1189_/A VGND VGND VPWR VPWR __dut__.__uuf__._1182_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1533__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__.__uuf__._2095__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1518_ __dut__.__uuf__._1509_/X __dut__.__uuf__._1505_/X __dut__._1168_/B
+ __dut__.__uuf__._1514_/X __dut__.__uuf__._1517_/X VGND VGND VPWR VPWR __dut__._1167_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1703_ __dut__._1719_/A1 __dut__._1701_/X __dut__._1702_/X VGND VGND VPWR
+ VPWR __dut__._1829_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1708__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1449_ __dut__.__uuf__._1449_/A VGND VGND VPWR VPWR __dut__.__uuf__._1449_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1669__A2 mp[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1634_ __dut__._1678_/A __dut__._1801_/Q VGND VGND VPWR VPWR __dut__._1634_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1565_ __dut__._1543_/Y mc[14] __dut__._1564_/X VGND VGND VPWR VPWR __dut__._1565_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1496_ rst VGND VGND VPWR VPWR __dut__._1496_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1443__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1357__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1109__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1618__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1303_ __dut__.__uuf__._1314_/A VGND VGND VPWR VPWR __dut__.__uuf__._1303_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1528__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1234_ __dut__.__uuf__._1249_/A VGND VGND VPWR VPWR __dut__.__uuf__._1234_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1165_ __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR __dut__.__uuf__._1165_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1096_ __dut__.__uuf__._1093_/X __dut__.__uuf__._1090_/X prod[57]
+ prod[58] __dut__.__uuf__._1085_/X VGND VGND VPWR VPWR __dut__._1383_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1350_ __dut__._1378_/A prod[40] VGND VGND VPWR VPWR __dut__._1350_/X sky130_fd_sc_hd__and2_4
X__dut__._1281_ __dut__._1281_/A1 __dut__._1281_/A2 __dut__._1280_/X VGND VGND VPWR
+ VPWR __dut__._1281_/X sky130_fd_sc_hd__a21o_4
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1587__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1998_ __dut__.__uuf__._1994_/Y __dut__.__uuf__._1995_/Y __dut__.__uuf__._1276_/X
+ __dut__.__uuf__._1997_/X VGND VGND VPWR VPWR __dut__.__uuf__._1999_/A sky130_fd_sc_hd__a211o_4
X_160_ _193_/B VGND VGND VPWR VPWR _172_/B sky130_fd_sc_hd__buf_2
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0996_ __dut__._1378_/A __dut__._1914_/Q VGND VGND VPWR VPWR __dut__._0996_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1438__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1617_ __dut__._1543_/Y mc[26] __dut__._1616_/X VGND VGND VPWR VPWR __dut__._1617_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1548_ __dut__._1788_/A __dut__._1791_/Q VGND VGND VPWR VPWR __dut__._1548_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1479_ rst VGND VGND VPWR VPWR __dut__._1479_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1872__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_289_ _314_/CLK _289_/D VGND VGND VPWR VPWR _289_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1348__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_171_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1708__A __dut__._1617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1921_ __dut__.__uuf__._1917_/Y __dut__.__uuf__._1918_/Y __dut__.__uuf__._1886_/X
+ __dut__.__uuf__._1920_/X VGND VGND VPWR VPWR __dut__.__uuf__._1922_/A sky130_fd_sc_hd__a211o_4
XFILLER_52_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1852_ __dut__._1072_/B VGND VGND VPWR VPWR __dut__.__uuf__._1852_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1569__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1783_ __dut__.__uuf__._1804_/A __dut__.__uuf__._1783_/B __dut__.__uuf__._1783_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1785_/B sky130_fd_sc_hd__or3_4
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1741__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1258__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2197_ __dut__.__uuf__._2200_/CLK __dut__._1383_/X __dut__.__uuf__._1095_/X
+ VGND VGND VPWR VPWR prod[57] sky130_fd_sc_hd__dfrtp_4
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1217_ __dut__.__uuf__._1212_/X __dut__.__uuf__._1209_/X prod[16]
+ prod[17] __dut__.__uuf__._1205_/X VGND VGND VPWR VPWR __dut__._1301_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_101_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1148_ __dut__.__uuf__._1159_/A VGND VGND VPWR VPWR __dut__.__uuf__._1148_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1402_ __dut__._1786_/A __dut__._1402_/B VGND VGND VPWR VPWR __dut__._1402_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_101_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1079_ __dut__.__uuf__._1075_/X __dut__.__uuf__._2003_/A prod[63]
+ __dut__._1132_/B __dut__.__uuf__._1069_/X VGND VGND VPWR VPWR __dut__._1395_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1333_ __dut__._1339_/A1 __dut__._1333_/A2 __dut__._1332_/X VGND VGND VPWR
+ VPWR __dut__._1333_/X sky130_fd_sc_hd__a21o_4
XFILLER_70_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1264_ __dut__._1786_/A __dut__._1264_/B VGND VGND VPWR VPWR __dut__._1264_/X
+ sky130_fd_sc_hd__and2_4
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1195_ __dut__._1779_/A1 __dut__._1195_/A2 __dut__._1194_/X VGND VGND VPWR
+ VPWR __dut__._1195_/X sky130_fd_sc_hd__a21o_4
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1895__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ _204_/Y _208_/X _211_/X _254_/Q _246_/Q VGND VGND VPWR VPWR tdo sky130_fd_sc_hd__a32o_4
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_143_ _295_/Q _296_/Q VGND VGND VPWR VPWR _220_/A sky130_fd_sc_hd__or2_4
XFILLER_51_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0979_ __dut__._0979_/A1 prod[21] __dut__._0978_/X VGND VGND VPWR VPWR __dut__._1906_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__.__uuf__._1083__B2 __dut__.__uuf__._1069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1723__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2120_ __dut__.__uuf__._2138_/CLK __dut__._1229_/X __dut__.__uuf__._1367_/X
+ VGND VGND VPWR VPWR __dut__._1230_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2051_ __dut__.__uuf__._2065_/CLK __dut__._1091_/X __dut__.__uuf__._1604_/X
+ VGND VGND VPWR VPWR __dut__._1092_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_96_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1541__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1904_ __dut__.__uuf__._1881_/X __dut__.__uuf__._1903_/B __dut__.__uuf__._1903_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1905_/C sky130_fd_sc_hd__o21ai_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1835_ __dut__.__uuf__._1835_/A VGND VGND VPWR VPWR __dut__._1069_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_52_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1766_ __dut__.__uuf__._1763_/Y __dut__.__uuf__._1764_/Y __dut__.__uuf__._1743_/X
+ __dut__.__uuf__._1770_/B VGND VGND VPWR VPWR __dut__.__uuf__._1766_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1697_ __dut__._1621_/X VGND VGND VPWR VPWR __dut__.__uuf__._1703_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._0902_ __dut__._1378_/A __dut__._1867_/Q VGND VGND VPWR VPWR __dut__._0902_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1882_ __dut__._1883_/CLK __dut__._1882_/D __dut__._1447_/Y VGND VGND VPWR
+ VPWR __dut__._1882_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1716__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_72_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1316_ __dut__._1316_/A prod[23] VGND VGND VPWR VPWR __dut__._1316_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2029__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1451__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1247_ __dut__._1787_/A1 __dut__._1247_/A2 __dut__._1246_/X VGND VGND VPWR
+ VPWR __dut__._1247_/X sky130_fd_sc_hd__a21o_4
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1178_ __dut__._1178_/A __dut__._1178_/B VGND VGND VPWR VPWR __dut__._1178_/X
+ sky130_fd_sc_hd__and2_4
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_126_ _256_/D _258_/D VGND VGND VPWR VPWR _127_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1910__CLK __dut__._1917_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1705__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_134_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1620_ __dut__.__uuf__._1624_/A VGND VGND VPWR VPWR __dut__.__uuf__._1620_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1551_ __dut__.__uuf__._1551_/A VGND VGND VPWR VPWR __dut__.__uuf__._1551_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1482_ __dut__.__uuf__._1486_/A VGND VGND VPWR VPWR __dut__.__uuf__._1482_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_89_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1536__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2103_ __dut__.__uuf__._2208_/CLK __dut__._1195_/X __dut__.__uuf__._1455_/X
+ VGND VGND VPWR VPWR __dut__._1196_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2034_ __dut__.__uuf__._2083_/CLK __dut__._1057_/X __dut__.__uuf__._1626_/X
+ VGND VGND VPWR VPWR __dut__._1058_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1101_ __dut__._1129_/A1 __dut__._1101_/A2 __dut__._1100_/X VGND VGND VPWR
+ VPWR __dut__._1101_/X sky130_fd_sc_hd__a21o_4
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1032_ __dut__._1078_/A __dut__._1032_/B VGND VGND VPWR VPWR __dut__._1032_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1818_ __dut__._1066_/B VGND VGND VPWR VPWR __dut__.__uuf__._1818_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1749_ __dut__.__uuf__._1749_/A __dut__.__uuf__._1749_/B __dut__.__uuf__._1749_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1751_/B sky130_fd_sc_hd__or3_4
X__dut__._1865_ __dut__._1915_/CLK __dut__._1865_/D __dut__._1464_/Y VGND VGND VPWR
+ VPWR __dut__._1865_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1446__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1796_ __dut__._1410_/B __dut__._1796_/D __dut__._1533_/Y VGND VGND VPWR
+ VPWR __dut__._1796_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_6_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__282__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1356__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1806__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1603_ __dut__.__uuf__._1605_/A VGND VGND VPWR VPWR __dut__.__uuf__._1603_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_30_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1534_ __dut__.__uuf__._1550_/A VGND VGND VPWR VPWR __dut__.__uuf__._1534_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1465_ __dut__.__uuf__._1465_/A VGND VGND VPWR VPWR __dut__.__uuf__._1465_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1650_ __dut__._1650_/A __dut__._1815_/Q VGND VGND VPWR VPWR __dut__._1650_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1396_ __dut__.__uuf__._1391_/X __dut__.__uuf__._1395_/X __dut__._1220_/B
+ __dut__.__uuf__._1391_/X VGND VGND VPWR VPWR __dut__._1219_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1581_ __dut__._1543_/Y mc[18] __dut__._1580_/X VGND VGND VPWR VPWR __dut__._1581_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1266__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2017_ __dut__.__uuf__._2049_/CLK __dut__._1023_/X __dut__.__uuf__._1646_/X
+ VGND VGND VPWR VPWR __dut__._1024_/B sky130_fd_sc_hd__dfrtp_4
Xclkbuf_4_6_0___dut__.__uuf__.__clk_source__ clkbuf_4_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2107_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_57_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1081__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_35_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1015_ __dut__._1129_/A1 __dut__._1015_/A2 __dut__._1014_/X VGND VGND VPWR
+ VPWR __dut__._1015_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1917_ __dut__._1917_/CLK __dut__._1917_/D __dut__._1412_/Y VGND VGND VPWR
+ VPWR __dut__._1917_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1848_ clkbuf_4_9_0_tck/X __dut__._1848_/D __dut__._1481_/Y VGND VGND VPWR
+ VPWR __dut__._1848_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._0895__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1779_ __dut__._1779_/A1 __dut__._1777_/X __dut__._1778_/X VGND VGND VPWR
+ VPWR __dut__._1848_/D sky130_fd_sc_hd__a21o_4
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1536__A __dut__.__uuf__._1536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_161 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._0882_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_150 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._0982_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_172 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1074_/A sky130_fd_sc_hd__buf_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_17 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0977_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_28 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0947_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_39 psn_inst_psn_buff_49/A VGND VGND VPWR VPWR __dut__._1301_/A1
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1250_ __dut__.__uuf__._1242_/X __dut__.__uuf__._1239_/X prod[5]
+ prod[6] __dut__.__uuf__._1249_/X VGND VGND VPWR VPWR __dut__._1279_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1181_ __dut__.__uuf__._1168_/X __dut__.__uuf__._1180_/X prod[29]
+ prod[30] __dut__.__uuf__._1175_/X VGND VGND VPWR VPWR __dut__._1327_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1086__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1063__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1517_ __dut__._1701_/X __dut__.__uuf__._1515_/X __dut__._1170_/B
+ __dut__.__uuf__._1516_/X VGND VGND VPWR VPWR __dut__.__uuf__._1517_/X sky130_fd_sc_hd__o22a_4
X__dut__._1702_ __dut__._1766_/A __dut__._1828_/Q VGND VGND VPWR VPWR __dut__._1702_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1448_ __dut__.__uuf__._1448_/A VGND VGND VPWR VPWR __dut__.__uuf__._1449_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_89_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1633_ __dut__._1543_/Y mc[2] __dut__._1632_/X VGND VGND VPWR VPWR __dut__._1633_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1379_ __dut__.__uuf__._1393_/A VGND VGND VPWR VPWR __dut__.__uuf__._1379_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1564_ __dut__._1788_/A __dut__._1795_/Q VGND VGND VPWR VPWR __dut__._1564_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1495_ rst VGND VGND VPWR VPWR __dut__._1495_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1724__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1634__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1045__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1302_ __dut__.__uuf__._1316_/A VGND VGND VPWR VPWR __dut__.__uuf__._1302_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1233_ __dut__.__uuf__._1233_/A VGND VGND VPWR VPWR __dut__.__uuf__._1233_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1164_ __dut__.__uuf__._1450_/A VGND VGND VPWR VPWR __dut__.__uuf__._1223_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1095_ __dut__.__uuf__._1099_/A VGND VGND VPWR VPWR __dut__.__uuf__._1095_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1280_ __dut__._1280_/A prod[5] VGND VGND VPWR VPWR __dut__._1280_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1997_ __dut__.__uuf__._1994_/Y __dut__.__uuf__._1995_/Y __dut__.__uuf__._1573_/A
+ __dut__.__uuf__._2001_/B VGND VGND VPWR VPWR __dut__.__uuf__._1997_/X sky130_fd_sc_hd__o22a_4
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0995_ __dut__._1327_/A1 prod[29] __dut__._0994_/X VGND VGND VPWR VPWR __dut__._1914_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1616_ __dut__._1788_/A __dut__._1808_/Q VGND VGND VPWR VPWR __dut__._1616_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1454__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1547_ __dut__._1647_/A1 __dut__._1545_/X __dut__._1546_/X VGND VGND VPWR
+ VPWR __dut__._1790_/D sky130_fd_sc_hd__a21o_4
XFILLER_92_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1478_ rst VGND VGND VPWR VPWR __dut__._1478_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1027__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__311__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_288_ _313_/CLK _288_/D VGND VGND VPWR VPWR _288_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_164_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1364__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1920_ __dut__.__uuf__._1917_/Y __dut__.__uuf__._1918_/Y __dut__.__uuf__._1908_/X
+ __dut__.__uuf__._1925_/B VGND VGND VPWR VPWR __dut__.__uuf__._1920_/X sky130_fd_sc_hd__o22a_4
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1851_ __dut__._1078_/B VGND VGND VPWR VPWR __dut__.__uuf__._1851_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1569__A2 mc[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1782_ __dut__.__uuf__._1774_/Y __dut__.__uuf__._1775_/Y __dut__.__uuf__._1774_/Y
+ __dut__.__uuf__._1775_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1783_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1539__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1741__A2 mp[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2196_ __dut__.__uuf__._2200_/CLK __dut__._1381_/X __dut__.__uuf__._1097_/X
+ VGND VGND VPWR VPWR prod[56] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1216_ __dut__.__uuf__._1218_/A VGND VGND VPWR VPWR __dut__.__uuf__._1216_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1147_ __dut__.__uuf__._1162_/A VGND VGND VPWR VPWR __dut__.__uuf__._1159_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1401_ __dut__._1787_/A1 __dut__._1401_/A2 __dut__._1400_/X VGND VGND VPWR
+ VPWR __dut__._1401_/X sky130_fd_sc_hd__a21o_4
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1332_ __dut__._1378_/A prod[31] VGND VGND VPWR VPWR __dut__._1332_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1257__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1078_ __dut__.__uuf__._1078_/A VGND VGND VPWR VPWR __dut__.__uuf__._2003_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1263_ __dut__._1787_/A1 __dut__._1263_/A2 __dut__._1262_/X VGND VGND VPWR
+ VPWR __dut__._1263_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1009__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1194_ __dut__._1194_/A __dut__._1194_/B VGND VGND VPWR VPWR __dut__._1194_/X
+ sky130_fd_sc_hd__and2_4
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ _211_/A _211_/B VGND VGND VPWR VPWR _211_/X sky130_fd_sc_hd__or2_4
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_142_ _296_/Q VGND VGND VPWR VPWR _142_/Y sky130_fd_sc_hd__inv_2
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1449__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0978_ __dut__._1404_/A __dut__._1905_/Q VGND VGND VPWR VPWR __dut__._0978_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1184__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1083__A2 __dut__.__uuf__._2003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1723__A2 __dut__._1721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2050_ __dut__.__uuf__._2065_/CLK __dut__._1089_/X __dut__.__uuf__._1605_/X
+ VGND VGND VPWR VPWR __dut__._1090_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1239__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1903_ __dut__.__uuf__._1914_/A __dut__.__uuf__._1903_/B __dut__.__uuf__._1903_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1905_/B sky130_fd_sc_hd__or3_4
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1834_ __dut__.__uuf__._1829_/Y __dut__.__uuf__._1830_/Y __dut__.__uuf__._1831_/X
+ __dut__.__uuf__._1833_/X VGND VGND VPWR VPWR __dut__.__uuf__._1835_/A sky130_fd_sc_hd__a211o_4
X__dut__.__uuf__._1765_ __dut__._1597_/X VGND VGND VPWR VPWR __dut__.__uuf__._1770_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1411__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2100__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._0901_ __dut__._1383_/A1 prod[47] __dut__._0900_/X VGND VGND VPWR VPWR __dut__._1867_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1696_ __dut__._1016_/B VGND VGND VPWR VPWR __dut__.__uuf__._1696_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1881_ __dut__._1883_/CLK __dut__._1881_/D __dut__._1448_/Y VGND VGND VPWR
+ VPWR __dut__._1881_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2179_ __dut__.__uuf__._2200_/CLK __dut__._1347_/X __dut__.__uuf__._1148_/X
+ VGND VGND VPWR VPWR prod[39] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1862__CLK __dut__._1917_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1315_ __dut__._1339_/A1 __dut__._1315_/A2 __dut__._1314_/X VGND VGND VPWR
+ VPWR __dut__._1315_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_65_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1732__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1246_ __dut__._1408_/A __dut__._1246_/B VGND VGND VPWR VPWR __dut__._1246_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1177_ __dut__._1647_/A1 __dut__._1177_/A2 __dut__._1176_/X VGND VGND VPWR
+ VPWR __dut__._1177_/X sky130_fd_sc_hd__a21o_4
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_125_ _237_/A _138_/B VGND VGND VPWR VPWR _125_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1705__A2 mp[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1641__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_127_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1550_ __dut__.__uuf__._1550_/A VGND VGND VPWR VPWR __dut__.__uuf__._1550_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1481_ __dut__.__uuf__._1466_/X __dut__.__uuf__._1462_/X __dut__._1184_/B
+ __dut__.__uuf__._1471_/X __dut__.__uuf__._1480_/X VGND VGND VPWR VPWR __dut__._1183_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_88_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2102_ __dut__.__uuf__._2208_/CLK __dut__._1193_/X __dut__.__uuf__._1458_/X
+ VGND VGND VPWR VPWR __dut__._1194_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2033_ __dut__.__uuf__._2083_/CLK __dut__._1055_/X __dut__.__uuf__._1627_/X
+ VGND VGND VPWR VPWR __dut__._1056_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1552__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1100_ __dut__._1100_/A __dut__._1100_/B VGND VGND VPWR VPWR __dut__._1100_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1031_ __dut__._1129_/A1 __dut__._1031_/A2 __dut__._1030_/X VGND VGND VPWR
+ VPWR __dut__._1031_/X sky130_fd_sc_hd__a21o_4
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1817_ __dut__.__uuf__._1828_/A __dut__.__uuf__._1817_/B __dut__.__uuf__._1817_/C
+ VGND VGND VPWR VPWR __dut__._1059_/A2 sky130_fd_sc_hd__and3_4
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1748_ __dut__.__uuf__._1741_/Y __dut__.__uuf__._1742_/Y __dut__.__uuf__._1741_/Y
+ __dut__.__uuf__._1742_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1749_/C sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1679_ __dut__.__uuf__._1673_/Y __dut__.__uuf__._1674_/Y __dut__.__uuf__._1673_/Y
+ __dut__.__uuf__._1674_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1680_/C sky130_fd_sc_hd__a2bb2o_4
X__dut__._1864_ __dut__._1915_/CLK __dut__._1864_/D __dut__._1465_/Y VGND VGND VPWR
+ VPWR __dut__._1864_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1795_ clkbuf_4_5_0_tck/X __dut__._1795_/D __dut__._1534_/Y VGND VGND VPWR
+ VPWR __dut__._1795_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1462__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2146__CLK __dut__.__uuf__._2164_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1623__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1229_ __dut__._1787_/A1 __dut__._1229_/A2 __dut__._1228_/X VGND VGND VPWR
+ VPWR __dut__._1229_/X sky130_fd_sc_hd__a21o_4
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1372__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1602_ __dut__.__uuf__._1605_/A VGND VGND VPWR VPWR __dut__.__uuf__._1602_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1533_ __dut__.__uuf__._1575_/A VGND VGND VPWR VPWR __dut__.__uuf__._1550_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2019__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1464_ __dut__.__uuf__._1443_/X __dut__.__uuf__._1462_/X __dut__._1192_/B
+ __dut__.__uuf__._1449_/X __dut__.__uuf__._1463_/X VGND VGND VPWR VPWR __dut__._1191_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_89_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1395_ __dut__.__uuf__._1394_/Y __dut__.__uuf__._1375_/X __dut__.__uuf__._1376_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1395_/X sky130_fd_sc_hd__o21a_4
X__dut__._1580_ __dut__._1788_/A __dut__._1799_/Q VGND VGND VPWR VPWR __dut__._1580_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_69_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2016_ __dut__.__uuf__._2049_/CLK __dut__._1021_/X __dut__.__uuf__._1647_/X
+ VGND VGND VPWR VPWR __dut__._1022_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1282__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1605__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1900__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1014_ __dut__._1128_/A __dut__._1014_/B VGND VGND VPWR VPWR __dut__._1014_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_28_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1440__A2 __dut__.__uuf__._1946_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1457__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1916_ __dut__._1917_/CLK __dut__._1916_/D __dut__._1413_/Y VGND VGND VPWR
+ VPWR __dut__._1916_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1847_ clkbuf_4_9_0_tck/X __dut__._1847_/D __dut__._1482_/Y VGND VGND VPWR
+ VPWR __dut__._1847_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1089__A __dut__.__uuf__._1450_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1778_ __dut__._1786_/A __dut__._1847_/Q VGND VGND VPWR VPWR __dut__._1778_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_162 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1346_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_151 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._0984_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_173 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1078_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_140 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1276_/A sky130_fd_sc_hd__buf_2
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_29 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._1283_/A1
+ sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_18 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0975_/A1
+ sky130_fd_sc_hd__buf_2
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1180_ __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR __dut__.__uuf__._1180_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1516_ __dut__.__uuf__._1720_/A VGND VGND VPWR VPWR __dut__.__uuf__._1516_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1701_ __dut__._1543_/Y mp[13] __dut__._1700_/X VGND VGND VPWR VPWR __dut__._1701_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1447_ __dut__.__uuf__._1465_/A VGND VGND VPWR VPWR __dut__.__uuf__._1447_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1632_ __dut__._1788_/A __dut__._1812_/Q VGND VGND VPWR VPWR __dut__._1632_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1378_ __dut__.__uuf__._1365_/X __dut__.__uuf__._1377_/X __dut__._1228_/B
+ __dut__.__uuf__._1365_/X VGND VGND VPWR VPWR __dut__._1227_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1563_ __dut__._1767_/A1 __dut__._1561_/X __dut__._1562_/X VGND VGND VPWR
+ VPWR __dut__._1794_/D sky130_fd_sc_hd__a21o_4
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__272__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1494_ rst VGND VGND VPWR VPWR __dut__._1494_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1740__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1301_ __dut__.__uuf__._1286_/X __dut__.__uuf__._1300_/X __dut__._1258_/B
+ __dut__.__uuf__._1286_/X VGND VGND VPWR VPWR __dut__._1257_/A2 sky130_fd_sc_hd__a2bb2o_4
XANTENNA__295__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1232_ __dut__.__uuf__._1227_/X __dut__.__uuf__._1223_/X prod[11]
+ prod[12] __dut__.__uuf__._1219_/X VGND VGND VPWR VPWR __dut__._1291_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1163_ __dut__.__uuf__._1174_/A VGND VGND VPWR VPWR __dut__.__uuf__._1163_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1094_ __dut__.__uuf__._1093_/X __dut__.__uuf__._1090_/X prod[58]
+ prod[59] __dut__.__uuf__._1085_/X VGND VGND VPWR VPWR __dut__._1385_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1544__B __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2207__CLK __dut__.__uuf__._2210_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1560__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1996_ __dut__._1545_/X VGND VGND VPWR VPWR __dut__.__uuf__._2001_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0904__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0994_ __dut__._1378_/A __dut__._1913_/Q VGND VGND VPWR VPWR __dut__._0994_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_2_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1615_ __dut__._1767_/A1 __dut__._1613_/X __dut__._1614_/X VGND VGND VPWR
+ VPWR __dut__._1807_/D sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_95_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1546_ tdi __dut__._1546_/B VGND VGND VPWR VPWR __dut__._1546_/X sky130_fd_sc_hd__and2_4
XFILLER_92_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1477_ rst VGND VGND VPWR VPWR __dut__._1477_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1470__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_287_ _314_/CLK _287_/D VGND VGND VPWR VPWR _287_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_psn_inst_psn_buff_157_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1380__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1850_ __dut__.__uuf__._1883_/A __dut__.__uuf__._1850_/B __dut__.__uuf__._1850_/C
+ VGND VGND VPWR VPWR __dut__._1071_/A2 sky130_fd_sc_hd__and3_4
XANTENNA___dut__.__uuf__._1086__B1 prod[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1781_ __dut__.__uuf__._1781_/A VGND VGND VPWR VPWR __dut__.__uuf__._1828_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2195_ __dut__.__uuf__._2200_/CLK __dut__._1379_/X __dut__.__uuf__._1099_/X
+ VGND VGND VPWR VPWR prod[55] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1215_ __dut__.__uuf__._1212_/X __dut__.__uuf__._1209_/X prod[17]
+ prod[18] __dut__.__uuf__._1205_/X VGND VGND VPWR VPWR __dut__._1303_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_101_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1146_ __dut__.__uuf__._1138_/X __dut__.__uuf__._1135_/X prod[40]
+ prod[41] __dut__.__uuf__._1145_/X VGND VGND VPWR VPWR __dut__._1349_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1400_ __dut__._1786_/A __dut__._1400_/B VGND VGND VPWR VPWR __dut__._1400_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_47_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1274__B prod[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1331_ __dut__._1331_/A1 __dut__._1331_/A2 __dut__._1330_/X VGND VGND VPWR
+ VPWR __dut__._1331_/X sky130_fd_sc_hd__a21o_4
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1077_ __dut__.__uuf__._1450_/A VGND VGND VPWR VPWR __dut__.__uuf__._1078_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1262_ __dut__._1786_/A __dut__._1262_/B VGND VGND VPWR VPWR __dut__._1262_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA__310__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1193_ __dut__._1193_/A1 __dut__._1193_/A2 __dut__._1192_/X VGND VGND VPWR
+ VPWR __dut__._1193_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1290__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1979_ __dut__.__uuf__._1936_/X __dut__.__uuf__._1978_/B __dut__.__uuf__._1978_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1980_/C sky130_fd_sc_hd__o21ai_4
XFILLER_23_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_210_ _209_/Y _210_/A2 _247_/Q _253_/Q VGND VGND VPWR VPWR _211_/B sky130_fd_sc_hd__o22a_4
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_141_ _295_/Q VGND VGND VPWR VPWR _239_/A sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1791__CLK __dut__._1410_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_10_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0977_ __dut__._0977_/A1 prod[20] __dut__._0976_/X VGND VGND VPWR VPWR __dut__._1905_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1465__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1529_ rst VGND VGND VPWR VPWR __dut__._1529_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1083__A3 prod[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1902_ __dut__.__uuf__._1896_/Y __dut__.__uuf__._1897_/Y __dut__.__uuf__._1896_/Y
+ __dut__.__uuf__._1897_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1903_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1833_ __dut__.__uuf__._1829_/Y __dut__.__uuf__._1830_/Y __dut__.__uuf__._1798_/X
+ __dut__.__uuf__._1838_/B VGND VGND VPWR VPWR __dut__.__uuf__._1833_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__._1411__A2 clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1764_ __dut__._1040_/B VGND VGND VPWR VPWR __dut__.__uuf__._1764_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1695_ __dut__._1022_/B VGND VGND VPWR VPWR __dut__.__uuf__._1695_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._0900_ __dut__._1378_/A __dut__._1866_/Q VGND VGND VPWR VPWR __dut__._0900_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1880_ __dut__._1883_/CLK __dut__._1880_/D __dut__._1449_/Y VGND VGND VPWR
+ VPWR __dut__._1880_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1175__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_tck clkbuf_4_9_0_tck/A VGND VGND VPWR VPWR clkbuf_4_9_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2178_ __dut__.__uuf__._2200_/CLK __dut__._1345_/X __dut__.__uuf__._1151_/X
+ VGND VGND VPWR VPWR prod[38] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1129_ __dut__.__uuf__._1124_/X __dut__.__uuf__._1121_/X prod[46]
+ prod[47] __dut__.__uuf__._1117_/X VGND VGND VPWR VPWR __dut__._1361_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_75_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1314_ __dut__._1314_/A prod[22] VGND VGND VPWR VPWR __dut__._1314_/X sky130_fd_sc_hd__and2_4
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1245_ __dut__._1787_/A1 __dut__._1245_/A2 __dut__._1244_/X VGND VGND VPWR
+ VPWR __dut__._1245_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_58_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1176_ __dut__._1176_/A __dut__._1176_/B VGND VGND VPWR VPWR __dut__._1176_/X
+ sky130_fd_sc_hd__and2_4
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_124_ _291_/Q VGND VGND VPWR VPWR _138_/B sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2075__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._0913__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1641__A2 mc[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1157__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1480_ __dut__._1737_/X __dut__.__uuf__._1472_/X __dut__._1186_/B
+ __dut__.__uuf__._1473_/X VGND VGND VPWR VPWR __dut__.__uuf__._1480_/X sky130_fd_sc_hd__o22a_4
XFILLER_88_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2101_ __dut__.__uuf__._2208_/CLK __dut__._1191_/X __dut__.__uuf__._1461_/X
+ VGND VGND VPWR VPWR __dut__._1192_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2032_ __dut__.__uuf__._2083_/CLK __dut__._1053_/X __dut__.__uuf__._1628_/X
+ VGND VGND VPWR VPWR __dut__._1054_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1030_ __dut__._1078_/A __dut__._1030_/B VGND VGND VPWR VPWR __dut__._1030_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1816_ __dut__.__uuf__._1771_/X __dut__.__uuf__._1815_/B __dut__.__uuf__._1815_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1817_/C sky130_fd_sc_hd__o21ai_4
XANTENNA___dut__.__uuf__._2098__CLK __dut__.__uuf__._2164_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1747_ __dut__.__uuf__._1747_/A VGND VGND VPWR VPWR __dut__._1037_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1678_ __dut__.__uuf__._1678_/A VGND VGND VPWR VPWR __dut__._1013_/A2
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._0912__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1863_ __dut__._1917_/CLK __dut__._1863_/D __dut__._1466_/Y VGND VGND VPWR
+ VPWR __dut__._1863_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1794_ clkbuf_4_5_0_tck/X __dut__._1794_/D __dut__._1535_/Y VGND VGND VPWR
+ VPWR __dut__._1794_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1623__A2 __dut__._1621_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1228_ __dut__._1786_/A __dut__._1228_/B VGND VGND VPWR VPWR __dut__._1228_/X
+ sky130_fd_sc_hd__and2_4
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1159_ __dut__._1159_/A1 __dut__._1159_/A2 __dut__._1158_/X VGND VGND VPWR
+ VPWR __dut__._1159_/X sky130_fd_sc_hd__a21o_4
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1139__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1601_ __dut__.__uuf__._1605_/A VGND VGND VPWR VPWR __dut__.__uuf__._1601_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1852__CLK __dut__._1410_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1532_ __dut__.__uuf__._1530_/X __dut__.__uuf__._1526_/X __dut__._1160_/B
+ __dut__.__uuf__._1514_/X __dut__.__uuf__._1531_/X VGND VGND VPWR VPWR __dut__._1159_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1463_ __dut__._1753_/X __dut__.__uuf__._1451_/X __dut__._1194_/B
+ __dut__.__uuf__._1452_/X VGND VGND VPWR VPWR __dut__.__uuf__._1463_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1394_ __dut__._1222_/B VGND VGND VPWR VPWR __dut__.__uuf__._1394_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._2015_ __dut__.__uuf__._2114_/CLK __dut__._1019_/X __dut__.__uuf__._1648_/X
+ VGND VGND VPWR VPWR __dut__._1020_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1605__A2 mc[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1013_ __dut__._1129_/A1 __dut__._1013_/A2 __dut__._1012_/X VGND VGND VPWR
+ VPWR __dut__._1013_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1369__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1915_ __dut__._1915_/CLK __dut__._1915_/D __dut__._1414_/Y VGND VGND VPWR
+ VPWR __dut__._1915_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1738__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1846_ __dut__._1902_/CLK __dut__._1846_/D __dut__._1483_/Y VGND VGND VPWR
+ VPWR __dut__._1846_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._2113__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1777_ __dut__._1543_/Y mp[30] __dut__._1776_/X VGND VGND VPWR VPWR __dut__._1777_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1473__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__305__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_130 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1192_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_163 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1378_/A sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_152 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1002_/A sky130_fd_sc_hd__buf_2
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_141 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._0944_/A sky130_fd_sc_hd__buf_2
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_174 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1128_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_19 psn_inst_psn_buff_9/A VGND VGND VPWR VPWR __dut__._0937_/A1
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1648__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1599__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1558__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1515_ __dut__.__uuf__._1536_/A VGND VGND VPWR VPWR __dut__.__uuf__._1515_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1700_ __dut__._1788_/A __dut__._1829_/Q VGND VGND VPWR VPWR __dut__._1700_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1446_ __dut__.__uuf__._1469_/A VGND VGND VPWR VPWR __dut__.__uuf__._1465_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1631_ __dut__._1647_/A1 __dut__._1629_/X __dut__._1630_/X VGND VGND VPWR
+ VPWR __dut__._1811_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1377_ __dut__.__uuf__._1374_/Y __dut__.__uuf__._1375_/X __dut__.__uuf__._1376_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1377_/X sky130_fd_sc_hd__o21a_4
X__dut__._1562_ __dut__._1766_/A __dut__._1793_/Q VGND VGND VPWR VPWR __dut__._1562_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1493_ rst VGND VGND VPWR VPWR __dut__._1493_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1898__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_40_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1468__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1829_ clkbuf_4_7_0_tck/X __dut__._1829_/D __dut__._1500_/Y VGND VGND VPWR
+ VPWR __dut__._1829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2009__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_102_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2159__CLK __dut__.__uuf__._2164_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1378__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1753__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1300_ __dut__.__uuf__._1294_/Y __dut__.__uuf__._1297_/X __dut__.__uuf__._1299_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1300_/X sky130_fd_sc_hd__o21a_4
XANTENNA__298__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1231_ __dut__.__uuf__._1233_/A VGND VGND VPWR VPWR __dut__.__uuf__._1231_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1162_ __dut__.__uuf__._1162_/A VGND VGND VPWR VPWR __dut__.__uuf__._1174_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_86_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1093_ __dut__.__uuf__._1138_/A VGND VGND VPWR VPWR __dut__.__uuf__._1093_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1995_ __dut__._1124_/B VGND VGND VPWR VPWR __dut__.__uuf__._1995_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_42_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1288__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0993_ __dut__._0993_/A1 prod[28] __dut__._0992_/X VGND VGND VPWR VPWR __dut__._1913_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1429_ __dut__._1208_/B VGND VGND VPWR VPWR __dut__.__uuf__._1429_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._0920__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1614_ __dut__._1766_/A __dut__._1806_/Q VGND VGND VPWR VPWR __dut__._1614_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1545_ mc[0] __dut__._1543_/Y __dut__._1544_/X VGND VGND VPWR VPWR __dut__._1545_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1476_ rst VGND VGND VPWR VPWR __dut__._1476_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_286_ _314_/CLK _286_/D VGND VGND VPWR VPWR _286_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1913__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1780_ __dut__.__uuf__._1780_/A VGND VGND VPWR VPWR __dut__._1049_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__262__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2194_ __dut__.__uuf__._2194_/CLK __dut__._1377_/X __dut__.__uuf__._1105_/X
+ VGND VGND VPWR VPWR prod[54] sky130_fd_sc_hd__dfrtp_4
XFILLER_87_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1214_ __dut__.__uuf__._1218_/A VGND VGND VPWR VPWR __dut__.__uuf__._1214_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1145_ __dut__.__uuf__._1175_/A VGND VGND VPWR VPWR __dut__.__uuf__._1145_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1330_ __dut__._1378_/A prod[30] VGND VGND VPWR VPWR __dut__._1330_/X sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1076_ __dut__.__uuf__._1438_/A VGND VGND VPWR VPWR __dut__.__uuf__._1450_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1261_ __dut__._1787_/A1 __dut__._1261_/A2 __dut__._1260_/X VGND VGND VPWR
+ VPWR __dut__._1261_/X sky130_fd_sc_hd__a21o_4
X__dut__._1192_ __dut__._1192_/A __dut__._1192_/B VGND VGND VPWR VPWR __dut__._1192_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_23_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1978_ __dut__.__uuf__._2001_/A __dut__.__uuf__._1978_/B __dut__.__uuf__._1978_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1980_/B sky130_fd_sc_hd__or3_4
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_140_ _140_/A VGND VGND VPWR VPWR _311_/D sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1717__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1746__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0976_ __dut__._1404_/A __dut__._1904_/Q VGND VGND VPWR VPWR __dut__._0976_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1528_ rst VGND VGND VPWR VPWR __dut__._1528_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1481__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1459_ rst VGND VGND VPWR VPWR __dut__._1459_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__285__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_269_ _314_/CLK _269_/D VGND VGND VPWR VPWR _269_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_6_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1656__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._0931__A2 prod[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1901_ __dut__.__uuf__._1901_/A VGND VGND VPWR VPWR __dut__._1093_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_37_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1832_ __dut__._1569_/X VGND VGND VPWR VPWR __dut__.__uuf__._1838_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1763_ __dut__._1046_/B VGND VGND VPWR VPWR __dut__.__uuf__._1763_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1694_ __dut__.__uuf__._1717_/A __dut__.__uuf__._1694_/B __dut__.__uuf__._1694_/C
+ VGND VGND VPWR VPWR __dut__._1015_/A2 sky130_fd_sc_hd__and3_4
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1566__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2177_ __dut__.__uuf__._2200_/CLK __dut__._1343_/X __dut__.__uuf__._1155_/X
+ VGND VGND VPWR VPWR prod[37] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1128_ __dut__.__uuf__._1130_/A VGND VGND VPWR VPWR __dut__.__uuf__._1128_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1313_ __dut__._1313_/A1 __dut__._1313_/A2 __dut__._1312_/X VGND VGND VPWR
+ VPWR __dut__._1313_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1059_ __dut__.__uuf__._1057_/Y __dut__.__uuf__._1058_/X __dut__.__uuf__._1054_/X
+ __dut__._1404_/B __dut__.__uuf__._1043_/X VGND VGND VPWR VPWR __dut__._1403_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1244_ __dut__._1786_/A __dut__._1244_/B VGND VGND VPWR VPWR __dut__._1244_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1175_ __dut__._1647_/A1 __dut__._1175_/A2 __dut__._1174_/X VGND VGND VPWR
+ VPWR __dut__._1175_/X sky130_fd_sc_hd__a21o_4
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_123_ _314_/Q VGND VGND VPWR VPWR _237_/A sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1476__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._0959_ __dut__._0961_/A1 prod[11] __dut__._0958_/X VGND VGND VPWR VPWR __dut__._1896_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_87_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1836__A __dut__.__uuf__._1946_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0___dut__.__uuf__.__clk_source__ clkbuf_2_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_46_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1386__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__300__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2100_ __dut__.__uuf__._2107_/CLK __dut__._1189_/X __dut__.__uuf__._1465_/X
+ VGND VGND VPWR VPWR __dut__._1190_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2031_ __dut__.__uuf__._2043_/CLK __dut__._1051_/X __dut__.__uuf__._1629_/X
+ VGND VGND VPWR VPWR __dut__._1052_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1093__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1815_ __dut__.__uuf__._1859_/A __dut__.__uuf__._1815_/B __dut__.__uuf__._1815_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1817_/B sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1746_ __dut__.__uuf__._1741_/Y __dut__.__uuf__._1742_/Y __dut__.__uuf__._1721_/X
+ __dut__.__uuf__._1745_/X VGND VGND VPWR VPWR __dut__.__uuf__._1747_/A sky130_fd_sc_hd__a211o_4
X__dut__.__uuf__._1677_ __dut__.__uuf__._1673_/Y __dut__.__uuf__._1674_/Y __dut__.__uuf__._1660_/X
+ __dut__.__uuf__._1676_/X VGND VGND VPWR VPWR __dut__.__uuf__._1678_/A sky130_fd_sc_hd__a211o_4
X__dut__._1862_ __dut__._1917_/CLK __dut__._1862_/D __dut__._1467_/Y VGND VGND VPWR
+ VPWR __dut__._1862_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1296__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1793_ __dut__._1410_/B __dut__._1793_/D __dut__._1536_/Y VGND VGND VPWR
+ VPWR __dut__._1793_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_psn_inst_psn_buff_70_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1227_ __dut__._1787_/A1 __dut__._1227_/A2 __dut__._1226_/X VGND VGND VPWR
+ VPWR __dut__._1227_/X sky130_fd_sc_hd__a21o_4
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1158_ __dut__._1766_/A __dut__._1158_/B VGND VGND VPWR VPWR __dut__._1158_/X
+ sky130_fd_sc_hd__and2_4
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1089_ __dut__._1129_/A1 __dut__._1089_/A2 __dut__._1088_/X VGND VGND VPWR
+ VPWR __dut__._1089_/X sky130_fd_sc_hd__a21o_4
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0_tck clkbuf_4_9_0_tck/A VGND VGND VPWR VPWR _290_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA_psn_inst_psn_buff_132_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1600_ __dut__.__uuf__._1606_/A VGND VGND VPWR VPWR __dut__.__uuf__._1605_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1531_ __dut__._1685_/X __dut__.__uuf__._1515_/X __dut__._1162_/B
+ __dut__.__uuf__._1516_/X VGND VGND VPWR VPWR __dut__.__uuf__._1531_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1462_ __dut__.__uuf__._1483_/A VGND VGND VPWR VPWR __dut__.__uuf__._1462_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._0889__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1393_ __dut__.__uuf__._1393_/A VGND VGND VPWR VPWR __dut__.__uuf__._1393_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2014_ __dut__.__uuf__._2114_/CLK __dut__._1017_/X __dut__.__uuf__._1650_/X
+ VGND VGND VPWR VPWR __dut__._1018_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1012_ __dut__._1128_/A __dut__._1012_/B VGND VGND VPWR VPWR __dut__._1012_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1729_ __dut__.__uuf__._1715_/X __dut__.__uuf__._1728_/B __dut__.__uuf__._1728_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1730_/C sky130_fd_sc_hd__o21ai_4
X__dut__._1914_ __dut__._1915_/CLK __dut__._1914_/D __dut__._1415_/Y VGND VGND VPWR
+ VPWR __dut__._1914_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1845_ clkbuf_4_5_0_tck/X __dut__._1845_/D __dut__._1484_/Y VGND VGND VPWR
+ VPWR __dut__._1845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1776_ __dut__._1788_/A __dut__._1848_/Q VGND VGND VPWR VPWR __dut__._1776_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1754__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_4_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xpsn_inst_psn_buff_120 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1590_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_164 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1542_/A sky130_fd_sc_hd__buf_4
Xpsn_inst_psn_buff_153 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1004_/A sky130_fd_sc_hd__buf_2
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpsn_inst_psn_buff_131 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1194_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_142 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1280_/A sky130_fd_sc_hd__buf_2
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_175 _236_/Y VGND VGND VPWR VPWR __dut__._1788_/A sky130_fd_sc_hd__buf_8
XFILLER_98_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1664__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1296__A __dut__.__uuf__._1720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1514_ __dut__.__uuf__._1535_/A VGND VGND VPWR VPWR __dut__.__uuf__._1514_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1445_ __dut__.__uuf__._1443_/X __dut__.__uuf__._1437_/X __dut__._1200_/B
+ __dut__.__uuf__._2004_/B __dut__.__uuf__._1444_/X VGND VGND VPWR VPWR __dut__._1199_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1630_ __dut__._1630_/A __dut__._1810_/Q VGND VGND VPWR VPWR __dut__._1630_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1376_ __dut__.__uuf__._1401_/A VGND VGND VPWR VPWR __dut__.__uuf__._1376_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_89_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1561_ __dut__._1543_/Y mc[13] __dut__._1560_/X VGND VGND VPWR VPWR __dut__._1561_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1574__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1492_ rst VGND VGND VPWR VPWR __dut__._1492_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._0918__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_33_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1211__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1828_ clkbuf_4_7_0_tck/X __dut__._1828_/D __dut__._1501_/Y VGND VGND VPWR
+ VPWR __dut__._1828_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1484__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1759_ __dut__._1759_/A1 __dut__._1757_/X __dut__._1758_/X VGND VGND VPWR
+ VPWR __dut__._1843_/D sky130_fd_sc_hd__a21o_4
XFILLER_49_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1842__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1753__A2 mp[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1230_ __dut__.__uuf__._1227_/X __dut__.__uuf__._1223_/X prod[12]
+ prod[13] __dut__.__uuf__._1219_/X VGND VGND VPWR VPWR __dut__._1293_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1394__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1161_ __dut__.__uuf__._1153_/X __dut__.__uuf__._1149_/X prod[35]
+ prod[36] __dut__.__uuf__._1160_/X VGND VGND VPWR VPWR __dut__._1339_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_86_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1092_ __dut__.__uuf__._1099_/A VGND VGND VPWR VPWR __dut__.__uuf__._1092_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1269__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1994_ __dut__._1134_/B VGND VGND VPWR VPWR __dut__.__uuf__._1994_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2103__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0992_ __dut__._1324_/A __dut__._1912_/Q VGND VGND VPWR VPWR __dut__._0992_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1428_ __dut__.__uuf__._1442_/A VGND VGND VPWR VPWR __dut__.__uuf__._1428_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1613_ __dut__._1543_/Y mc[25] __dut__._1612_/X VGND VGND VPWR VPWR __dut__._1613_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1359_ __dut__._1236_/B VGND VGND VPWR VPWR __dut__.__uuf__._1359_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1865__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1544_ __dut__._1790_/Q __dut__._1788_/A VGND VGND VPWR VPWR __dut__._1544_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1475_ rst VGND VGND VPWR VPWR __dut__._1475_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_2_0___dut__.__uuf__.__clk_source__ clkbuf_4_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2119_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_45_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1479__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_285_ _290_/CLK _285_/D VGND VGND VPWR VPWR _285_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1671__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1086__A2 __dut__.__uuf__._2003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1888__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1213_ __dut__.__uuf__._1212_/X __dut__.__uuf__._1209_/X prod[18]
+ prod[19] __dut__.__uuf__._1205_/X VGND VGND VPWR VPWR __dut__._1305_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._2193_ __dut__.__uuf__._2194_/CLK __dut__._1375_/X __dut__.__uuf__._1108_/X
+ VGND VGND VPWR VPWR prod[53] sky130_fd_sc_hd__dfrtp_4
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1144_ __dut__.__uuf__._1144_/A VGND VGND VPWR VPWR __dut__.__uuf__._1144_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1075_ __dut__.__uuf__._1138_/A VGND VGND VPWR VPWR __dut__.__uuf__._1075_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1260_ __dut__._1786_/A __dut__._1260_/B VGND VGND VPWR VPWR __dut__._1260_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_82_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1191_ __dut__._1193_/A1 __dut__._1191_/A2 __dut__._1190_/X VGND VGND VPWR
+ VPWR __dut__._1191_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1977_ __dut__.__uuf__._1971_/Y __dut__.__uuf__._1972_/Y __dut__.__uuf__._1971_/Y
+ __dut__.__uuf__._1972_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1978_/C sky130_fd_sc_hd__a2bb2o_4
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1717__A2 mp[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0975_ __dut__._0975_/A1 prod[19] __dut__._0974_/X VGND VGND VPWR VPWR __dut__._1904_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_tck clkbuf_0_tck/X VGND VGND VPWR VPWR clkbuf_2_3_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1762__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1527_ rst VGND VGND VPWR VPWR __dut__._1527_/Y sky130_fd_sc_hd__inv_2
X__dut__._1458_ rst VGND VGND VPWR VPWR __dut__._1458_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1653__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1389_ __dut__._1389_/A1 __dut__._1389_/A2 __dut__._1388_/X VGND VGND VPWR
+ VPWR __dut__._1389_/X sky130_fd_sc_hd__a21o_4
XFILLER_14_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_268_ _313_/CLK _268_/D VGND VGND VPWR VPWR _268_/Q sky130_fd_sc_hd__dfxtp_4
X_199_ _199_/A VGND VGND VPWR VPWR _199_/X sky130_fd_sc_hd__buf_2
XFILLER_96_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_162_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1672__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1900_ __dut__.__uuf__._1896_/Y __dut__.__uuf__._1897_/Y __dut__.__uuf__._1886_/X
+ __dut__.__uuf__._1899_/X VGND VGND VPWR VPWR __dut__.__uuf__._1901_/A sky130_fd_sc_hd__a211o_4
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1831_ __dut__.__uuf__._1941_/A VGND VGND VPWR VPWR __dut__.__uuf__._1831_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1762_ __dut__.__uuf__._1773_/A __dut__.__uuf__._1762_/B __dut__.__uuf__._1762_/C
+ VGND VGND VPWR VPWR __dut__._1039_/A2 sky130_fd_sc_hd__and3_4
X__dut__.__uuf__._1693_ __dut__.__uuf__._1573_/X __dut__.__uuf__._1692_/B __dut__.__uuf__._1692_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1694_/C sky130_fd_sc_hd__o21ai_4
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2176_ __dut__.__uuf__._2200_/CLK __dut__._1341_/X __dut__.__uuf__._1157_/X
+ VGND VGND VPWR VPWR prod[36] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1127_ __dut__.__uuf__._1124_/X __dut__.__uuf__._1121_/X prod[47]
+ prod[48] __dut__.__uuf__._1117_/X VGND VGND VPWR VPWR __dut__._1363_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1582__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1058_ __dut__._1404_/B __dut__.__uuf__._1058_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1058_/X sky130_fd_sc_hd__or2_4
X__dut__._1312_ __dut__._1404_/A prod[21] VGND VGND VPWR VPWR __dut__._1312_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1635__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1243_ __dut__._1787_/A1 __dut__._1243_/A2 __dut__._1242_/X VGND VGND VPWR
+ VPWR __dut__._1243_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._1942__A __dut__._1765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._0926__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1174_ __dut__._1174_/A __dut__._1174_/B VGND VGND VPWR VPWR __dut__._1174_/X
+ sky130_fd_sc_hd__and2_4
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_122_ _291_/Q VGND VGND VPWR VPWR _231_/A sky130_fd_sc_hd__buf_2
X__dut__._0958_ __dut__._1770_/A __dut__._1895_/Q VGND VGND VPWR VPWR __dut__._0958_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0889_ __dut__._1383_/A1 prod[41] __dut__._0888_/X VGND VGND VPWR VPWR __dut__._1861_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_87_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1492__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2030_ __dut__.__uuf__._2083_/CLK __dut__._1049_/X __dut__.__uuf__._1630_/X
+ VGND VGND VPWR VPWR __dut__._1050_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1617__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1814_ __dut__.__uuf__._1807_/Y __dut__.__uuf__._1808_/Y __dut__.__uuf__._1807_/Y
+ __dut__.__uuf__._1808_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1815_/C sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1745_ __dut__.__uuf__._1741_/Y __dut__.__uuf__._1742_/Y __dut__.__uuf__._1743_/X
+ __dut__.__uuf__._1749_/B VGND VGND VPWR VPWR __dut__.__uuf__._1745_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1676_ __dut__.__uuf__._1673_/Y __dut__.__uuf__._1674_/Y __dut__.__uuf__._2001_/A
+ __dut__.__uuf__._1680_/B VGND VGND VPWR VPWR __dut__.__uuf__._1676_/X sky130_fd_sc_hd__o22a_4
X__dut__._1861_ __dut__._1917_/CLK __dut__._1861_/D __dut__._1468_/Y VGND VGND VPWR
+ VPWR __dut__._1861_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1792_ __dut__._1410_/B __dut__._1792_/D __dut__._1537_/Y VGND VGND VPWR
+ VPWR __dut__._1792_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__275__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2159_ __dut__.__uuf__._2164_/CLK __dut__._1307_/X __dut__.__uuf__._1208_/X
+ VGND VGND VPWR VPWR prod[19] sky130_fd_sc_hd__dfrtp_4
XFILLER_28_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_63_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1226_ __dut__._1786_/A __dut__._1226_/B VGND VGND VPWR VPWR __dut__._1226_/X
+ sky130_fd_sc_hd__and2_4
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1157_ __dut__._1767_/A1 __dut__._1157_/A2 __dut__._1156_/X VGND VGND VPWR
+ VPWR __dut__._1157_/X sky130_fd_sc_hd__a21o_4
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1088_ __dut__._1094_/A __dut__._1088_/B VGND VGND VPWR VPWR __dut__._1088_/X
+ sky130_fd_sc_hd__and2_4
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1487__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2008__A __dut__.__uuf__._2008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_125_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1530_ __dut__.__uuf__._1551_/A VGND VGND VPWR VPWR __dut__.__uuf__._1530_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1461_ __dut__.__uuf__._1465_/A VGND VGND VPWR VPWR __dut__.__uuf__._1461_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1392_ __dut__.__uuf__._1380_/X __dut__.__uuf__._1390_/X __dut__._1222_/B
+ __dut__.__uuf__._1391_/X VGND VGND VPWR VPWR __dut__._1221_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2013_ __dut__.__uuf__._2114_/CLK __dut__._1015_/X __dut__.__uuf__._1651_/X
+ VGND VGND VPWR VPWR __dut__._1016_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_69_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1011_ __dut__._1129_/A1 __dut__._1011_/A2 __dut__._1010_/X VGND VGND VPWR
+ VPWR __dut__._1011_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1728_ __dut__.__uuf__._1749_/A __dut__.__uuf__._1728_/B __dut__.__uuf__._1728_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1730_/B sky130_fd_sc_hd__or3_4
X__dut__._1913_ __dut__._1915_/CLK __dut__._1913_/D __dut__._1416_/Y VGND VGND VPWR
+ VPWR __dut__._1913_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1659_ __dut__._1128_/B VGND VGND VPWR VPWR __dut__.__uuf__._1659_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1844_ __dut__._1899_/CLK __dut__._1844_/D __dut__._1485_/Y VGND VGND VPWR
+ VPWR __dut__._1844_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1775_ __dut__._1779_/A1 __dut__._1773_/X __dut__._1774_/X VGND VGND VPWR
+ VPWR __dut__._1847_/D sky130_fd_sc_hd__a21o_4
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1770__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpsn_inst_psn_buff_110 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1044_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_121 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1130_/A sky130_fd_sc_hd__buf_2
XFILLER_44_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1209_ __dut__._1787_/A1 __dut__._1209_/A2 __dut__._1208_/X VGND VGND VPWR
+ VPWR __dut__._1209_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_154 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1338_/A sky130_fd_sc_hd__buf_2
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_132 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1198_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_143 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._0970_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_165 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1324_/A sky130_fd_sc_hd__buf_2
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__314__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1680__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1513_ __dut__.__uuf__._1529_/A VGND VGND VPWR VPWR __dut__.__uuf__._1513_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1444_ __dut__._1773_/X __dut__.__uuf__._1946_/A __dut__._1202_/B
+ __dut__.__uuf__._1425_/X VGND VGND VPWR VPWR __dut__.__uuf__._1444_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1375_ __dut__.__uuf__._1400_/A VGND VGND VPWR VPWR __dut__.__uuf__._1375_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_89_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1560_ __dut__._1788_/A __dut__._1794_/Q VGND VGND VPWR VPWR __dut__._1560_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2032__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1487__A __dut__.__uuf__._1551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1491_ rst VGND VGND VPWR VPWR __dut__._1491_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1794__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_26_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_tck clkbuf_4_7_0_tck/A VGND VGND VPWR VPWR clkbuf_4_7_0_tck/X sky130_fd_sc_hd__clkbuf_1
X__dut__._1827_ clkbuf_4_7_0_tck/X __dut__._1827_/D __dut__._1502_/Y VGND VGND VPWR
+ VPWR __dut__._1827_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1758_ __dut__._1770_/A __dut__._1842_/Q VGND VGND VPWR VPWR __dut__._1758_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1689_ __dut__._1543_/Y mp[10] __dut__._1688_/X VGND VGND VPWR VPWR __dut__._1689_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_95_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1394__B prod[62] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1160_ __dut__.__uuf__._1175_/A VGND VGND VPWR VPWR __dut__.__uuf__._1160_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1100__A __dut__.__uuf__._1100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1091_ __dut__.__uuf__._1075_/X __dut__.__uuf__._1090_/X prod[59]
+ prod[60] __dut__.__uuf__._1085_/X VGND VGND VPWR VPWR __dut__._1387_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1993_ __dut__._1130_/B __dut__.__uuf__._1991_/X __dut__._1129_/A2
+ VGND VGND VPWR VPWR __dut__._1127_/A2 sky130_fd_sc_hd__a21boi_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0991_ __dut__._0991_/A1 prod[27] __dut__._0990_/X VGND VGND VPWR VPWR __dut__._1912_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1427_ __dut__.__uuf__._1416_/X __dut__.__uuf__._1426_/X __dut__._1208_/B
+ __dut__.__uuf__._1416_/X VGND VGND VPWR VPWR __dut__._1207_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1612_ __dut__._1788_/A __dut__._1807_/Q VGND VGND VPWR VPWR __dut__._1612_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1358_ __dut__.__uuf__._1367_/A VGND VGND VPWR VPWR __dut__.__uuf__._1358_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1543_ __dut__._1788_/A VGND VGND VPWR VPWR __dut__._1543_/Y sky130_fd_sc_hd__inv_8
X__dut__.__uuf__._1289_ __dut__._1262_/B VGND VGND VPWR VPWR __dut__.__uuf__._1289_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1474_ rst VGND VGND VPWR VPWR __dut__._1474_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_284_ _290_/CLK _284_/D VGND VGND VPWR VPWR _284_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2078__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1495__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1086__A3 prod[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0___dut__.__uuf__.__clk_source__ clkbuf_3_6_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2164_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_9_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1212_ __dut__.__uuf__._1212_/A VGND VGND VPWR VPWR __dut__.__uuf__._1212_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2192_ __dut__.__uuf__._2194_/CLK __dut__._1373_/X __dut__.__uuf__._1111_/X
+ VGND VGND VPWR VPWR prod[52] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1143_ __dut__.__uuf__._1138_/X __dut__.__uuf__._1135_/X prod[41]
+ prod[42] __dut__.__uuf__._1131_/X VGND VGND VPWR VPWR __dut__._1351_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1074_ __dut__.__uuf__._1551_/A VGND VGND VPWR VPWR __dut__.__uuf__._1138_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1111__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1190_ __dut__._1190_/A __dut__._1190_/B VGND VGND VPWR VPWR __dut__._1190_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1976_ __dut__.__uuf__._1976_/A VGND VGND VPWR VPWR __dut__._1121_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1832__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0974_ __dut__._0974_/A __dut__._1903_/Q VGND VGND VPWR VPWR __dut__._0974_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_93_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1526_ rst VGND VGND VPWR VPWR __dut__._1526_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1457_ rst VGND VGND VPWR VPWR __dut__._1457_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1653__A2 mp[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1388_ __dut__._1542_/A prod[59] VGND VGND VPWR VPWR __dut__._1388_/X sky130_fd_sc_hd__and2_4
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1169__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_267_ _313_/CLK _267_/D VGND VGND VPWR VPWR _267_/Q sky130_fd_sc_hd__dfxtp_4
X_198_ _199_/A VGND VGND VPWR VPWR _198_/X sky130_fd_sc_hd__buf_2
XFILLER_6_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_155_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1830_ __dut__._1064_/B VGND VGND VPWR VPWR __dut__.__uuf__._1830_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1761_ __dut__.__uuf__._1715_/X __dut__.__uuf__._1760_/B __dut__.__uuf__._1760_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1762_/C sky130_fd_sc_hd__o21ai_4
XANTENNA___dut__._1855__CLK __dut__._1919_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1692_ __dut__.__uuf__._1692_/A __dut__.__uuf__._1692_/B __dut__.__uuf__._1692_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1694_/B sky130_fd_sc_hd__or3_4
XANTENNA___dut__._0907__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2175_ __dut__.__uuf__._2200_/CLK __dut__._1339_/X __dut__.__uuf__._1159_/X
+ VGND VGND VPWR VPWR prod[35] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1126_ __dut__.__uuf__._1130_/A VGND VGND VPWR VPWR __dut__.__uuf__._1126_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_87_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1057_ __dut__.__uuf__._1057_/A VGND VGND VPWR VPWR __dut__.__uuf__._1057_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1311_ __dut__._1311_/A1 __dut__._1311_/A2 __dut__._1310_/X VGND VGND VPWR
+ VPWR __dut__._1311_/X sky130_fd_sc_hd__a21o_4
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1242_ __dut__._1786_/A __dut__._1242_/B VGND VGND VPWR VPWR __dut__._1242_/X
+ sky130_fd_sc_hd__and2_4
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1399__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1173_ __dut__._1647_/A1 __dut__._1173_/A2 __dut__._1172_/X VGND VGND VPWR
+ VPWR __dut__._1173_/X sky130_fd_sc_hd__a21o_4
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1959_ __dut__.__uuf__._1936_/X __dut__.__uuf__._1958_/B __dut__.__uuf__._1958_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1960_/C sky130_fd_sc_hd__o21ai_4
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_121_ _310_/Q VGND VGND VPWR VPWR _121_/Y sky130_fd_sc_hd__inv_2
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1571__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2116__CLK __dut__.__uuf__._2119_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._0957_ __dut__._0961_/A1 prod[10] __dut__._0956_/X VGND VGND VPWR VPWR __dut__._1895_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0888_ __dut__._1378_/A __dut__._1860_/Q VGND VGND VPWR VPWR __dut__._0888_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_78_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1509_ rst VGND VGND VPWR VPWR __dut__._1509_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1878__CLK __dut__._1919_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1617__A2 mc[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_tck clkbuf_0_tck/X VGND VGND VPWR VPWR clkbuf_2_1_0_tck/A sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1813_ __dut__.__uuf__._1868_/A VGND VGND VPWR VPWR __dut__.__uuf__._1859_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1744_ __dut__._1605_/X VGND VGND VPWR VPWR __dut__.__uuf__._1749_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1675_ __dut__._1629_/X VGND VGND VPWR VPWR __dut__.__uuf__._1680_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2139__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1860_ __dut__._1917_/CLK __dut__._1860_/D __dut__._1469_/Y VGND VGND VPWR
+ VPWR __dut__._1860_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1791_ __dut__._1410_/B __dut__._1791_/D __dut__._1538_/Y VGND VGND VPWR
+ VPWR __dut__._1791_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1553__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2158_ __dut__.__uuf__._2164_/CLK __dut__._1305_/X __dut__.__uuf__._1211_/X
+ VGND VGND VPWR VPWR prod[18] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1109_ __dut__.__uuf__._1138_/A VGND VGND VPWR VPWR __dut__.__uuf__._1109_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2089_ __dut__.__uuf__._2097_/CLK __dut__._1167_/X __dut__.__uuf__._1513_/X
+ VGND VGND VPWR VPWR __dut__._1168_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1953__A __dut__._1721_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_56_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1225_ __dut__._1787_/A1 __dut__._1225_/A2 __dut__._1224_/X VGND VGND VPWR
+ VPWR __dut__._1225_/X sky130_fd_sc_hd__a21o_4
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1156_ __dut__._1766_/A __dut__._1156_/B VGND VGND VPWR VPWR __dut__._1156_/X
+ sky130_fd_sc_hd__and2_4
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1087_ __dut__._1129_/A1 __dut__._1087_/A2 __dut__._1086_/X VGND VGND VPWR
+ VPWR __dut__._1087_/X sky130_fd_sc_hd__a21o_4
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1768__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_118_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1678__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1783__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1460_ __dut__.__uuf__._1443_/X __dut__.__uuf__._1437_/X __dut__._1194_/B
+ __dut__.__uuf__._1449_/X __dut__.__uuf__._1459_/X VGND VGND VPWR VPWR __dut__._1193_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__.__uuf__._1103__A __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1391_ __dut__.__uuf__._1416_/A VGND VGND VPWR VPWR __dut__.__uuf__._1391_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2012_ __dut__.__uuf__._2114_/CLK __dut__._1013_/X __dut__.__uuf__._1652_/X
+ VGND VGND VPWR VPWR __dut__._1014_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1010_ __dut__._1128_/A __dut__._1010_/B VGND VGND VPWR VPWR __dut__._1010_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1588__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1727_ __dut__.__uuf__._1718_/Y __dut__.__uuf__._1719_/Y __dut__.__uuf__._1718_/Y
+ __dut__.__uuf__._1719_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1728_/C sky130_fd_sc_hd__a2bb2o_4
X__dut__._1912_ __dut__._1915_/CLK __dut__._1912_/D __dut__._1417_/Y VGND VGND VPWR
+ VPWR __dut__._1912_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1658_ __dut__._1010_/B VGND VGND VPWR VPWR __dut__.__uuf__._1658_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1843_ __dut__._1899_/CLK __dut__._1843_/D __dut__._1486_/Y VGND VGND VPWR
+ VPWR __dut__._1843_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1589_ __dut__.__uuf__._1593_/A VGND VGND VPWR VPWR __dut__.__uuf__._1589_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1774_ __dut__._1774_/A __dut__._1846_/Q VGND VGND VPWR VPWR __dut__._1774_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpsn_inst_psn_buff_100 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1102_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_111 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1042_/A sky130_fd_sc_hd__buf_2
X__dut__._1208_ __dut__._1786_/A __dut__._1208_/B VGND VGND VPWR VPWR __dut__._1208_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_155 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1344_/A sky130_fd_sc_hd__buf_2
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_122 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1546_/B sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_133 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1774_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_144 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1770_/A sky130_fd_sc_hd__buf_4
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1139_ __dut__._1647_/A1 __dut__._1139_/A2 __dut__._1138_/X VGND VGND VPWR
+ VPWR __dut__._1139_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1498__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_166 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1308_/A sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1916__CLK __dut__._1917_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1765__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1512_ __dut__.__uuf__._1575_/A VGND VGND VPWR VPWR __dut__.__uuf__._1529_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1443_ __dut__.__uuf__._1466_/A VGND VGND VPWR VPWR __dut__.__uuf__._1443_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1374_ __dut__._1230_/B VGND VGND VPWR VPWR __dut__.__uuf__._1374_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1490_ rst VGND VGND VPWR VPWR __dut__._1490_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_psn_inst_psn_buff_19_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._0950__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1826_ clkbuf_4_7_0_tck/X __dut__._1826_/D __dut__._1503_/Y VGND VGND VPWR
+ VPWR __dut__._1826_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1757_ __dut__._1543_/Y mp[26] __dut__._1756_/X VGND VGND VPWR VPWR __dut__._1757_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1688_ __dut__._1788_/A __dut__._1826_/Q VGND VGND VPWR VPWR __dut__._1688_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_95_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1090_ __dut__.__uuf__._1149_/A VGND VGND VPWR VPWR __dut__.__uuf__._1090_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1992_ __dut__._1130_/B __dut__.__uuf__._1991_/X __dut__.__uuf__._1781_/A
+ VGND VGND VPWR VPWR __dut__._1129_/A2 sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._1729__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._0990_ __dut__._1324_/A __dut__._1911_/Q VGND VGND VPWR VPWR __dut__._0990_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1426_ __dut__.__uuf__._1424_/Y __dut__.__uuf__._1425_/X __dut__.__uuf__._1324_/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._1426_/X sky130_fd_sc_hd__o21a_4
X__dut__._1611_ __dut__._1767_/A1 __dut__._1609_/X __dut__._1610_/X VGND VGND VPWR
+ VPWR __dut__._1806_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1357_ __dut__.__uuf__._1354_/X __dut__.__uuf__._1356_/X __dut__._1236_/B
+ __dut__.__uuf__._1354_/X VGND VGND VPWR VPWR __dut__._1235_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1542_ __dut__._1542_/A VGND VGND VPWR VPWR __dut__._1542_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1288_ __dut__.__uuf__._1288_/A VGND VGND VPWR VPWR __dut__.__uuf__._1288_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1473_ rst VGND VGND VPWR VPWR __dut__._1473_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_283_ _290_/CLK _283_/D VGND VGND VPWR VPWR _283_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1776__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._0943__A2 prod[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1809_ clkbuf_4_7_0_tck/X __dut__._1809_/D __dut__._1520_/Y VGND VGND VPWR
+ VPWR __dut__._1809_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_100_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2022__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_9_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1686__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1211_ __dut__.__uuf__._1218_/A VGND VGND VPWR VPWR __dut__.__uuf__._1211_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2191_ __dut__.__uuf__._2194_/CLK __dut__._1371_/X __dut__.__uuf__._1113_/X
+ VGND VGND VPWR VPWR prod[51] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1142_ __dut__.__uuf__._1144_/A VGND VGND VPWR VPWR __dut__.__uuf__._1142_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1073_ __dut__.__uuf__._1226_/A VGND VGND VPWR VPWR __dut__.__uuf__._1551_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_6_0_tck clkbuf_4_7_0_tck/A VGND VGND VPWR VPWR clkbuf_4_6_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1975_ __dut__.__uuf__._1971_/Y __dut__.__uuf__._1972_/Y __dut__.__uuf__._1941_/X
+ __dut__.__uuf__._1974_/X VGND VGND VPWR VPWR __dut__.__uuf__._1976_/A sky130_fd_sc_hd__a211o_4
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._0925__A2 prod[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1596__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0973_ __dut__._1319_/A1 prod[18] __dut__._0972_/X VGND VGND VPWR VPWR __dut__._1903_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1409_ __dut__.__uuf__._1418_/A VGND VGND VPWR VPWR __dut__.__uuf__._1409_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1525_ rst VGND VGND VPWR VPWR __dut__._1525_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1456_ rst VGND VGND VPWR VPWR __dut__._1456_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1387_ __dut__._1387_/A1 __dut__._1387_/A2 __dut__._1386_/X VGND VGND VPWR
+ VPWR __dut__._1387_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2045__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_266_ _314_/CLK _266_/D VGND VGND VPWR VPWR _266_/Q sky130_fd_sc_hd__dfxtp_4
X_197_ _199_/A VGND VGND VPWR VPWR _197_/X sky130_fd_sc_hd__buf_2
XFILLER_96_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_psn_inst_psn_buff_148_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1760_ __dut__.__uuf__._1804_/A __dut__.__uuf__._1760_/B __dut__.__uuf__._1760_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1762_/B sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1691_ __dut__.__uuf__._1683_/Y __dut__.__uuf__._1684_/Y __dut__.__uuf__._1683_/Y
+ __dut__.__uuf__._1684_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1692_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2174_ __dut__.__uuf__._2194_/CLK __dut__._1337_/X __dut__.__uuf__._1163_/X
+ VGND VGND VPWR VPWR prod[34] sky130_fd_sc_hd__dfrtp_4
XFILLER_101_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1125_ __dut__.__uuf__._1124_/X __dut__.__uuf__._1121_/X prod[48]
+ prod[49] __dut__.__uuf__._1117_/X VGND VGND VPWR VPWR __dut__._1365_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1310_ __dut__._1404_/A prod[20] VGND VGND VPWR VPWR __dut__._1310_/X sky130_fd_sc_hd__and2_4
XFILLER_28_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2068__CLK __dut__.__uuf__._2119_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1056_ __dut__.__uuf__._1063_/A VGND VGND VPWR VPWR __dut__.__uuf__._1056_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_28_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1241_ __dut__._1787_/A1 __dut__._1241_/A2 __dut__._1240_/X VGND VGND VPWR
+ VPWR __dut__._1241_/X sky130_fd_sc_hd__a21o_4
XFILLER_83_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__291__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1172_ __dut__._1174_/A __dut__._1172_/B VGND VGND VPWR VPWR __dut__._1172_/X
+ sky130_fd_sc_hd__and2_4
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1958_ __dut__.__uuf__._1968_/A __dut__.__uuf__._1958_/B __dut__.__uuf__._1958_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1960_/B sky130_fd_sc_hd__or3_4
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1889_ __dut__.__uuf__._1884_/Y __dut__.__uuf__._1885_/Y __dut__.__uuf__._1886_/X
+ __dut__.__uuf__._1888_/X VGND VGND VPWR VPWR __dut__.__uuf__._1890_/A sky130_fd_sc_hd__a211o_4
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0956_ __dut__._1770_/A __dut__._1894_/Q VGND VGND VPWR VPWR __dut__._0956_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._0887_ __dut__._1349_/A1 prod[40] __dut__._0886_/X VGND VGND VPWR VPWR __dut__._1860_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_78_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1087__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1508_ rst VGND VGND VPWR VPWR __dut__._1508_/Y sky130_fd_sc_hd__inv_2
XANTENNA__308__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1439_ rst VGND VGND VPWR VPWR __dut__._1439_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_249_ _200_/X _313_/Q VGND VGND VPWR VPWR _249_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1011__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2210__CLK __dut__.__uuf__._2210_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_84_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1812_ __dut__.__uuf__._1812_/A VGND VGND VPWR VPWR __dut__._1061_/A2
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1204__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1743_ __dut__.__uuf__._1923_/A VGND VGND VPWR VPWR __dut__.__uuf__._1743_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1674_ __dut__._1008_/B VGND VGND VPWR VPWR __dut__.__uuf__._1674_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1553__A2 mc[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1790_ _194_/A __dut__._1790_/D __dut__._1539_/Y VGND VGND VPWR VPWR __dut__._1790_/Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2157_ __dut__.__uuf__._2169_/CLK __dut__._1303_/X __dut__.__uuf__._1214_/X
+ VGND VGND VPWR VPWR prod[17] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1108_ __dut__.__uuf__._1115_/A VGND VGND VPWR VPWR __dut__.__uuf__._1108_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2088_ __dut__.__uuf__._2097_/CLK __dut__._1165_/X __dut__.__uuf__._1519_/X
+ VGND VGND VPWR VPWR __dut__._1166_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1039_ __dut__.__uuf__._1438_/A VGND VGND VPWR VPWR __dut__.__uuf__._1295_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1224_ __dut__._1786_/A __dut__._1224_/B VGND VGND VPWR VPWR __dut__._1224_/X
+ sky130_fd_sc_hd__and2_4
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1114__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_49_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1155_ __dut__._1155_/A1 __dut__._1155_/A2 __dut__._1154_/X VGND VGND VPWR
+ VPWR __dut__._1155_/X sky130_fd_sc_hd__a21o_4
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1086_ __dut__._1678_/A __dut__._1086_/B VGND VGND VPWR VPWR __dut__._1086_/X
+ sky130_fd_sc_hd__and2_4
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1241__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1784__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0939_ __dut__._0939_/A1 prod[1] __dut__._0938_/X VGND VGND VPWR VPWR __dut__._1886_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_78_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1845__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1390_ __dut__.__uuf__._1389_/Y __dut__.__uuf__._1375_/X __dut__.__uuf__._1376_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1390_/X sky130_fd_sc_hd__o21a_4
XANTENNA___dut__._1694__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._2011_ __dut__.__uuf__._2114_/CLK __dut__._1011_/X __dut__.__uuf__._1653_/X
+ VGND VGND VPWR VPWR __dut__._1012_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_97_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2106__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1223__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1726_ __dut__.__uuf__._1781_/A VGND VGND VPWR VPWR __dut__.__uuf__._1773_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_21_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1911_ __dut__._1915_/CLK __dut__._1911_/D __dut__._1418_/Y VGND VGND VPWR
+ VPWR __dut__._1911_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1657_ __dut__.__uuf__._1657_/A VGND VGND VPWR VPWR done sky130_fd_sc_hd__buf_2
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1588_ __dut__.__uuf__._1606_/A VGND VGND VPWR VPWR __dut__.__uuf__._1593_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1842_ __dut__._1899_/CLK __dut__._1842_/D __dut__._1487_/Y VGND VGND VPWR
+ VPWR __dut__._1842_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1868__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1773_ __dut__._1543_/Y mp[29] __dut__._1772_/X VGND VGND VPWR VPWR __dut__._1773_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2209_ __dut__.__uuf__._2210_/CLK __dut__._1407_/X __dut__.__uuf__._1063_/A
+ VGND VGND VPWR VPWR __dut__._1408_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._0948__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_101 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1100_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_112 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1626_/A sky130_fd_sc_hd__buf_2
X__dut__._1207_ __dut__._1787_/A1 __dut__._1207_/A2 __dut__._1206_/X VGND VGND VPWR
+ VPWR __dut__._1207_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_145 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1304_/A sky130_fd_sc_hd__buf_2
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1138_ __dut__._1138_/A __dut__._1138_/B VGND VGND VPWR VPWR __dut__._1138_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_123 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1176_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_134 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1200_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_156 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1340_/A sky130_fd_sc_hd__buf_2
XFILLER_12_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_167 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1404_/A sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1765__A2 mc[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1069_ __dut__._1071_/A1 __dut__._1069_/A2 __dut__._1068_/X VGND VGND VPWR
+ VPWR __dut__._1069_/X sky130_fd_sc_hd__a21o_4
XFILLER_8_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_130_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1205__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1511_ __dut__.__uuf__._1509_/X __dut__.__uuf__._1505_/X __dut__._1170_/B
+ __dut__.__uuf__._1493_/X __dut__.__uuf__._1510_/X VGND VGND VPWR VPWR __dut__._1169_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1442_ __dut__.__uuf__._1442_/A VGND VGND VPWR VPWR __dut__.__uuf__._1442_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1373_ __dut__.__uuf__._1393_/A VGND VGND VPWR VPWR __dut__.__uuf__._1373_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1709_ __dut__.__uuf__._1706_/Y __dut__.__uuf__._1707_/Y __dut__.__uuf__._1686_/X
+ __dut__.__uuf__._1713_/B VGND VGND VPWR VPWR __dut__.__uuf__._1709_/X sky130_fd_sc_hd__o22a_4
X__dut__._1825_ clkbuf_4_7_0_tck/X __dut__._1825_/D __dut__._1504_/Y VGND VGND VPWR
+ VPWR __dut__._1825_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1756_ __dut__._1788_/A __dut__._1843_/Q VGND VGND VPWR VPWR __dut__._1756_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_95_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1687_ __dut__._1719_/A1 __dut__._1685_/X __dut__._1686_/X VGND VGND VPWR
+ VPWR __dut__._1825_/D sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_2_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1683__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1991_ __dut__._1140_/B __dut__._1641_/X VGND VGND VPWR VPWR __dut__.__uuf__._1991_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1729__A2 mp[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1212__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1425_ __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR __dut__.__uuf__._1425_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1610_ __dut__._1766_/A __dut__._1805_/Q VGND VGND VPWR VPWR __dut__._1610_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1356_ __dut__.__uuf__._1355_/Y __dut__.__uuf__._1349_/X __dut__.__uuf__._1350_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1356_/X sky130_fd_sc_hd__o21a_4
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1541_ rst VGND VGND VPWR VPWR __dut__._1541_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1287_ __dut__.__uuf__._1274_/X __dut__.__uuf__._1285_/X __dut__._1262_/B
+ __dut__.__uuf__._1286_/X VGND VGND VPWR VPWR __dut__._1261_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1472_ rst VGND VGND VPWR VPWR __dut__._1472_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1665__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1906__CLK __dut__._1919_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1122__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_282_ _290_/CLK _282_/D VGND VGND VPWR VPWR _282_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_psn_inst_psn_buff_31_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1808_ clkbuf_4_5_0_tck/X __dut__._1808_/D __dut__._1521_/Y VGND VGND VPWR
+ VPWR __dut__._1808_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1739_ __dut__._1739_/A1 __dut__._1737_/X __dut__._1738_/X VGND VGND VPWR
+ VPWR __dut__._1838_/D sky130_fd_sc_hd__a21o_4
XFILLER_76_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2190_ __dut__.__uuf__._2194_/CLK __dut__._1369_/X __dut__.__uuf__._1115_/X
+ VGND VGND VPWR VPWR prod[50] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1210_ __dut__.__uuf__._1198_/X __dut__.__uuf__._1209_/X prod[19]
+ prod[20] __dut__.__uuf__._1205_/X VGND VGND VPWR VPWR __dut__._1307_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1141_ __dut__.__uuf__._1138_/X __dut__.__uuf__._1135_/X prod[42]
+ prod[43] __dut__.__uuf__._1131_/X VGND VGND VPWR VPWR __dut__._1353_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1072_ __dut__.__uuf__._1084_/A VGND VGND VPWR VPWR __dut__.__uuf__._1072_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1647__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1974_ __dut__.__uuf__._1971_/Y __dut__.__uuf__._1972_/Y __dut__.__uuf__._1573_/A
+ __dut__.__uuf__._1978_/B VGND VGND VPWR VPWR __dut__.__uuf__._1974_/X sky130_fd_sc_hd__o22a_4
XFILLER_35_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0972_ __dut__._1308_/A __dut__._1902_/Q VGND VGND VPWR VPWR __dut__._0972_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__278__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1408_ __dut__.__uuf__._1405_/X __dut__.__uuf__._1407_/X __dut__._1216_/B
+ __dut__.__uuf__._1405_/X VGND VGND VPWR VPWR __dut__._1215_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1339_ __dut__.__uuf__._1338_/Y __dut__.__uuf__._1323_/X __dut__.__uuf__._1324_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1339_/X sky130_fd_sc_hd__o21a_4
X__dut__._1524_ rst VGND VGND VPWR VPWR __dut__._1524_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_79_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1455_ rst VGND VGND VPWR VPWR __dut__._1455_/Y sky130_fd_sc_hd__inv_2
XANTENNA__306__SET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1386_ __dut__._1542_/A prod[58] VGND VGND VPWR VPWR __dut__._1386_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._0956__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_265_ _313_/CLK _265_/D VGND VGND VPWR VPWR _265_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_196_ _199_/A VGND VGND VPWR VPWR _196_/X sky130_fd_sc_hd__buf_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1629__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._0866__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1690_ __dut__.__uuf__._1690_/A VGND VGND VPWR VPWR __dut__._1017_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_99_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2173_ __dut__.__uuf__._2194_/CLK __dut__._1335_/X __dut__.__uuf__._1167_/X
+ VGND VGND VPWR VPWR prod[33] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1124_ __dut__.__uuf__._1138_/A VGND VGND VPWR VPWR __dut__.__uuf__._1124_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1055_ __dut__.__uuf__._1052_/Y __dut__.__uuf__._1053_/X __dut__.__uuf__._1054_/X
+ __dut__._1406_/B __dut__.__uuf__._1043_/X VGND VGND VPWR VPWR __dut__._1405_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1240_ __dut__._1786_/A __dut__._1240_/B VGND VGND VPWR VPWR __dut__._1240_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1171_ __dut__._1647_/A1 __dut__._1171_/A2 __dut__._1170_/X VGND VGND VPWR
+ VPWR __dut__._1171_/X sky130_fd_sc_hd__a21o_4
XFILLER_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1957_ __dut__.__uuf__._1951_/Y __dut__.__uuf__._1952_/Y __dut__.__uuf__._1951_/Y
+ __dut__.__uuf__._1952_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1958_/C sky130_fd_sc_hd__a2bb2o_4
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1888_ __dut__.__uuf__._1884_/Y __dut__.__uuf__._1885_/Y __dut__.__uuf__._1853_/X
+ __dut__.__uuf__._1893_/B VGND VGND VPWR VPWR __dut__.__uuf__._1888_/X sky130_fd_sc_hd__o22a_4
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1400__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0955_ __dut__._0961_/A1 prod[9] __dut__._0954_/X VGND VGND VPWR VPWR __dut__._1894_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0886_ __dut__._1378_/A __dut__._1859_/Q VGND VGND VPWR VPWR __dut__._0886_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2012__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1507_ rst VGND VGND VPWR VPWR __dut__._1507_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1438_ rst VGND VGND VPWR VPWR __dut__._1438_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__.__uuf__._2162__CLK __dut__.__uuf__._2164_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1369_ __dut__._1383_/A1 __dut__._1369_/A2 __dut__._1368_/X VGND VGND VPWR
+ VPWR __dut__._1369_/X sky130_fd_sc_hd__a21o_4
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_248_ _201_/X _312_/Q VGND VGND VPWR VPWR _248_/Q sky130_fd_sc_hd__dfxtp_4
X_179_ _273_/Q _182_/B VGND VGND VPWR VPWR _272_/D sky130_fd_sc_hd__and2_4
Xclkbuf_4_5_0_tck clkbuf_4_5_0_tck/A VGND VGND VPWR VPWR clkbuf_4_5_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_160_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1811_ __dut__.__uuf__._1807_/Y __dut__.__uuf__._1808_/Y __dut__.__uuf__._1776_/X
+ __dut__.__uuf__._1810_/X VGND VGND VPWR VPWR __dut__.__uuf__._1812_/A sky130_fd_sc_hd__a211o_4
X__dut__.__uuf__._1742_ __dut__._1032_/B VGND VGND VPWR VPWR __dut__.__uuf__._1742_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_33_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1673_ __dut__._1014_/B VGND VGND VPWR VPWR __dut__.__uuf__._1673_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1220__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2035__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2156_ __dut__.__uuf__._2169_/CLK __dut__._1301_/X __dut__.__uuf__._1216_/X
+ VGND VGND VPWR VPWR prod[16] sky130_fd_sc_hd__dfrtp_4
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1107_ __dut__.__uuf__._1093_/X __dut__.__uuf__._1106_/X prod[54]
+ prod[55] __dut__.__uuf__._1100_/X VGND VGND VPWR VPWR __dut__._1377_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_75_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2087_ __dut__.__uuf__._2097_/CLK __dut__._1163_/X __dut__.__uuf__._1522_/X
+ VGND VGND VPWR VPWR __dut__._1164_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1038_ __dut__._1136_/B __dut__._1138_/B VGND VGND VPWR VPWR __dut__.__uuf__._1438_/A
+ sky130_fd_sc_hd__or2_4
X__dut__._1223_ __dut__._1787_/A1 __dut__._1223_/A2 __dut__._1222_/X VGND VGND VPWR
+ VPWR __dut__._1223_/X sky130_fd_sc_hd__a21o_4
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1797__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1154_ __dut__._1766_/A __dut__._1154_/B VGND VGND VPWR VPWR __dut__._1154_/X
+ sky130_fd_sc_hd__and2_4
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1085_ __dut__._1129_/A1 __dut__._1085_/A2 __dut__._1084_/X VGND VGND VPWR
+ VPWR __dut__._1085_/X sky130_fd_sc_hd__a21o_4
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1697__A __dut__._1621_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0938_ __dut__._1404_/A __dut__._1885_/Q VGND VGND VPWR VPWR __dut__._0938_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_79_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._0869_ __dut__._1543_/Y mc[8] __dut__._0868_/X VGND VGND VPWR VPWR __dut__._0869_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._2010_ __dut__.__uuf__._2119_/CLK __dut__._1009_/X __dut__.__uuf__._1654_/X
+ VGND VGND VPWR VPWR __dut__._1010_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_38_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1725_ __dut__.__uuf__._1725_/A VGND VGND VPWR VPWR __dut__._1029_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_33_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1910_ __dut__._1917_/CLK __dut__._1910_/D __dut__._1419_/Y VGND VGND VPWR
+ VPWR __dut__._1910_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1656_ __dut__.__uuf__._2005_/A __dut__._1138_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1657_/A sky130_fd_sc_hd__and2_4
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1587_ __dut__.__uuf__._1587_/A VGND VGND VPWR VPWR __dut__.__uuf__._1587_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1841_ __dut__._1899_/CLK __dut__._1841_/D __dut__._1488_/Y VGND VGND VPWR
+ VPWR __dut__._1841_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1772_ __dut__._1788_/A __dut__._1847_/Q VGND VGND VPWR VPWR __dut__._1772_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2208_ __dut__.__uuf__._2208_/CLK __dut__._1405_/X __dut__.__uuf__._1051_/X
+ VGND VGND VPWR VPWR __dut__._1406_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2139_ __dut__.__uuf__._2208_/CLK __dut__._1267_/X __dut__.__uuf__._1266_/X
+ VGND VGND VPWR VPWR __dut__._1268_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_61_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpsn_inst_psn_buff_102 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1098_/A sky130_fd_sc_hd__buf_2
X__dut__._1206_ __dut__._1786_/A __dut__._1206_/B VGND VGND VPWR VPWR __dut__._1206_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpsn_inst_psn_buff_146 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1302_/A sky130_fd_sc_hd__buf_2
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_113 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1630_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_124 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1174_/A sky130_fd_sc_hd__buf_2
X__dut__._1137_ __dut__._1779_/A1 __dut__._1137_/A2 __dut__._1136_/X VGND VGND VPWR
+ VPWR __dut__._1137_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_135 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1272_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_157 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._0876_/A sky130_fd_sc_hd__buf_2
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_168 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1786_/A sky130_fd_sc_hd__buf_8
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1068_ __dut__._1074_/A __dut__._1068_/B VGND VGND VPWR VPWR __dut__._1068_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_98_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._0874__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_123_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1510_ __dut__._1705_/X __dut__.__uuf__._1494_/X __dut__._1172_/B
+ __dut__.__uuf__._1495_/X VGND VGND VPWR VPWR __dut__.__uuf__._1510_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1441_ __dut__.__uuf__._1257_/X __dut__.__uuf__._1437_/X __dut__._1202_/B
+ __dut__.__uuf__._2004_/B __dut__.__uuf__._1440_/X VGND VGND VPWR VPWR __dut__._1201_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1372_ __dut__.__uuf__._1469_/A VGND VGND VPWR VPWR __dut__.__uuf__._1393_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1141__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1264__B1 prod[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1708_ __dut__._1617_/X VGND VGND VPWR VPWR __dut__.__uuf__._1713_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1835__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1639_ __dut__.__uuf__._1642_/A VGND VGND VPWR VPWR __dut__.__uuf__._1639_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1824_ clkbuf_4_7_0_tck/X __dut__._1824_/D __dut__._1505_/Y VGND VGND VPWR
+ VPWR __dut__._1824_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1755_ __dut__._1759_/A1 __dut__._1753_/X __dut__._1754_/X VGND VGND VPWR
+ VPWR __dut__._1842_/D sky130_fd_sc_hd__a21o_4
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1686_ __dut__._1766_/A __dut__._1824_/Q VGND VGND VPWR VPWR __dut__._1686_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1371__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1123__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1990_ __dut__.__uuf__._1990_/A __dut__.__uuf__._1990_/B __dut__.__uuf__._1990_/C
+ VGND VGND VPWR VPWR __dut__._1123_/A2 sky130_fd_sc_hd__and3_4
XFILLER_23_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1424_ __dut__._1210_/B VGND VGND VPWR VPWR __dut__.__uuf__._1424_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1355_ __dut__._1238_/B VGND VGND VPWR VPWR __dut__.__uuf__._1355_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1540_ rst VGND VGND VPWR VPWR __dut__._1540_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1286_ __dut__.__uuf__._1314_/A VGND VGND VPWR VPWR __dut__.__uuf__._1286_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1471_ rst VGND VGND VPWR VPWR __dut__._1471_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1665__A2 mp[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_281_ _290_/CLK _281_/D VGND VGND VPWR VPWR _281_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_psn_inst_psn_buff_24_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2119__CLK __dut__.__uuf__._2119_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1353__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1807_ clkbuf_4_5_0_tck/X __dut__._1807_/D __dut__._1522_/Y VGND VGND VPWR
+ VPWR __dut__._1807_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1105__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1738_ __dut__._1770_/A __dut__._1837_/Q VGND VGND VPWR VPWR __dut__._1738_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1669_ __dut__._1543_/Y mp[6] __dut__._1668_/X VGND VGND VPWR VPWR __dut__._1669_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._0919__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1140_ __dut__.__uuf__._1144_/A VGND VGND VPWR VPWR __dut__.__uuf__._1140_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1071_ __dut__._1398_/B __dut__.__uuf__._1069_/X __dut__.__uuf__._1029_/B
+ __dut__.__uuf__._1070_/X VGND VGND VPWR VPWR __dut__._1397_/A2 sky130_fd_sc_hd__o22a_4
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1973_ __dut__._1633_/X VGND VGND VPWR VPWR __dut__.__uuf__._1978_/B
+ sky130_fd_sc_hd__inv_2
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1583__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0971_ __dut__._1319_/A1 prod[17] __dut__._0970_/X VGND VGND VPWR VPWR __dut__._1902_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1407_ __dut__.__uuf__._1406_/Y __dut__.__uuf__._1400_/X __dut__.__uuf__._1401_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1407_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1338_ __dut__._1244_/B VGND VGND VPWR VPWR __dut__.__uuf__._1338_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1523_ rst VGND VGND VPWR VPWR __dut__._1523_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1269_ __dut__.__uuf__._1535_/A VGND VGND VPWR VPWR __dut__.__uuf__._2004_/B
+ sky130_fd_sc_hd__buf_2
X__dut__._1454_ rst VGND VGND VPWR VPWR __dut__._1454_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1385_ __dut__._1385_/A1 __dut__._1385_/A2 __dut__._1384_/X VGND VGND VPWR
+ VPWR __dut__._1385_/X sky130_fd_sc_hd__a21o_4
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_264_ _313_/CLK _264_/D VGND VGND VPWR VPWR _264_/Q sky130_fd_sc_hd__dfxtp_4
X_195_ _203_/A VGND VGND VPWR VPWR _199_/A sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._2091__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1629__A2 mc[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1565__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__312__SET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2172_ __dut__.__uuf__._2194_/CLK __dut__._1333_/X __dut__.__uuf__._1170_/X
+ VGND VGND VPWR VPWR prod[32] sky130_fd_sc_hd__dfrtp_4
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1123_ __dut__.__uuf__._1130_/A VGND VGND VPWR VPWR __dut__.__uuf__._1123_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1218__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1054_ __dut__.__uuf__._1100_/A VGND VGND VPWR VPWR __dut__.__uuf__._1054_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_28_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1170_ __dut__._1174_/A __dut__._1170_/B VGND VGND VPWR VPWR __dut__._1170_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1956_ __dut__.__uuf__._1956_/A VGND VGND VPWR VPWR __dut__._1113_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1887_ __dut__._1549_/X VGND VGND VPWR VPWR __dut__.__uuf__._1893_/B
+ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_1_1_0_tck_A clkbuf_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0954_ __dut__._1770_/A __dut__._1893_/Q VGND VGND VPWR VPWR __dut__._0954_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._0885_ __dut__._1349_/A1 prod[39] __dut__._0884_/X VGND VGND VPWR VPWR __dut__._1859_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_91_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1506_ rst VGND VGND VPWR VPWR __dut__._1506_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1437_ rst VGND VGND VPWR VPWR __dut__._1437_/Y sky130_fd_sc_hd__inv_2
X__dut__._1368_ __dut__._1378_/A prod[49] VGND VGND VPWR VPWR __dut__._1368_/X sky130_fd_sc_hd__and2_4
X__dut__._1299_ __dut__._1299_/A1 __dut__._1299_/A2 __dut__._1298_/X VGND VGND VPWR
+ VPWR __dut__._1299_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1919__CLK __dut__._1919_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1547__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_247_ _202_/X _311_/Q VGND VGND VPWR VPWR _247_/Q sky130_fd_sc_hd__dfxtp_4
X_178_ _274_/Q _182_/B VGND VGND VPWR VPWR _273_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1038__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_153_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1810_ __dut__.__uuf__._1807_/Y __dut__.__uuf__._1808_/Y __dut__.__uuf__._1798_/X
+ __dut__.__uuf__._1815_/B VGND VGND VPWR VPWR __dut__.__uuf__._1810_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1741_ __dut__._1038_/B VGND VGND VPWR VPWR __dut__.__uuf__._1741_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1501__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1672_ __dut__.__uuf__._1717_/A __dut__.__uuf__._1672_/B __dut__.__uuf__._1672_/C
+ VGND VGND VPWR VPWR __dut__._1007_/A2 sky130_fd_sc_hd__and3_4
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2155_ __dut__.__uuf__._2169_/CLK __dut__._1299_/X __dut__.__uuf__._1218_/X
+ VGND VGND VPWR VPWR prod[15] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1106_ __dut__.__uuf__._1149_/A VGND VGND VPWR VPWR __dut__.__uuf__._1106_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_75_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2086_ __dut__.__uuf__._2097_/CLK __dut__._1161_/X __dut__.__uuf__._1525_/X
+ VGND VGND VPWR VPWR __dut__._1162_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1037_ __dut__._0936_/B __dut__.__uuf__._1037_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1037_/X sky130_fd_sc_hd__or2_4
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1222_ __dut__._1786_/A __dut__._1222_/B VGND VGND VPWR VPWR __dut__._1222_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1153_ __dut__._1153_/A1 __dut__._1153_/A2 __dut__._1152_/X VGND VGND VPWR
+ VPWR __dut__._1153_/X sky130_fd_sc_hd__a21o_4
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1939_ __dut__._1110_/B VGND VGND VPWR VPWR __dut__.__uuf__._1939_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_12_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1084_ __dut__._1084_/A __dut__._1084_/B VGND VGND VPWR VPWR __dut__._1084_/X
+ sky130_fd_sc_hd__and2_4
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1777__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._0937_ __dut__._0937_/A1 prod[0] __dut__._0936_/X VGND VGND VPWR VPWR __dut__._1885_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0868_ __dut__._1788_/A __dut__._1853_/Q VGND VGND VPWR VPWR __dut__._0868_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1701__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1891__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1724_ __dut__.__uuf__._1718_/Y __dut__.__uuf__._1719_/Y __dut__.__uuf__._1721_/X
+ __dut__.__uuf__._1723_/X VGND VGND VPWR VPWR __dut__.__uuf__._1725_/A sky130_fd_sc_hd__a211o_4
X__dut__.__uuf__._1655_ __dut__.__uuf__._2008_/A VGND VGND VPWR VPWR __dut__.__uuf__._1655_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1586_ __dut__.__uuf__._1587_/A VGND VGND VPWR VPWR __dut__.__uuf__._1586_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1840_ __dut__._1899_/CLK __dut__._1840_/D __dut__._1489_/Y VGND VGND VPWR
+ VPWR __dut__._1840_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1771_ __dut__._1771_/A1 __dut__._1769_/X __dut__._1770_/X VGND VGND VPWR
+ VPWR __dut__._1846_/D sky130_fd_sc_hd__a21o_4
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2207_ __dut__.__uuf__._2210_/CLK __dut__._1403_/X __dut__.__uuf__._1056_/X
+ VGND VGND VPWR VPWR __dut__._1404_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._2138_ __dut__.__uuf__._2138_/CLK __dut__._1265_/X __dut__.__uuf__._1273_/X
+ VGND VGND VPWR VPWR __dut__._1266_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_75_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2069_ __dut__.__uuf__._2119_/CLK __dut__._1127_/X __dut__.__uuf__._1583_/X
+ VGND VGND VPWR VPWR __dut__._1128_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA__245__A1 tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_103 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1094_/A sky130_fd_sc_hd__buf_2
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_54_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1205_ __dut__._1787_/A1 __dut__._1205_/A2 __dut__._1204_/X VGND VGND VPWR
+ VPWR __dut__._1205_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_4_4_0_tck clkbuf_4_5_0_tck/A VGND VGND VPWR VPWR __dut__._1410_/B sky130_fd_sc_hd__clkbuf_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_114 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1638_/A sky130_fd_sc_hd__buf_2
X__dut__._1136_ __dut__._1786_/A __dut__._1136_/B VGND VGND VPWR VPWR __dut__._1136_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_125 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1178_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_136 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1270_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_158 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1408_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_147 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1318_/A sky130_fd_sc_hd__buf_2
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xpsn_inst_psn_buff_169 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1274_/A sky130_fd_sc_hd__buf_2
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1067_ __dut__._1071_/A1 __dut__._1067_/A2 __dut__._1066_/X VGND VGND VPWR
+ VPWR __dut__._1067_/X sky130_fd_sc_hd__a21o_4
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_116_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._0890__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1440_ __dut__._1777_/X __dut__.__uuf__._1946_/A __dut__._1204_/B
+ __dut__.__uuf__._1425_/X VGND VGND VPWR VPWR __dut__.__uuf__._1440_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1371_ __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR __dut__.__uuf__._1469_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_2_0_0_tck_A clkbuf_2_1_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0___dut__.__uuf__.__clk_source__ clkbuf_4_7_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2097_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1226__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1707_ __dut__._1020_/B VGND VGND VPWR VPWR __dut__.__uuf__._1707_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1638_ __dut__.__uuf__._1642_/A VGND VGND VPWR VPWR __dut__.__uuf__._1638_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1823_ clkbuf_4_5_0_tck/X __dut__._1823_/D __dut__._1506_/Y VGND VGND VPWR
+ VPWR __dut__._1823_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1569_ __dut__.__uuf__._1569_/A VGND VGND VPWR VPWR __dut__.__uuf__._1569_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1754_ __dut__._1770_/A __dut__._1841_/Q VGND VGND VPWR VPWR __dut__._1754_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1685_ __dut__._1543_/Y mp[9] __dut__._1684_/X VGND VGND VPWR VPWR __dut__._1685_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1136__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._0891__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2048__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1119_ __dut__._1129_/A1 __dut__._1119_/A2 __dut__._1118_/X VGND VGND VPWR
+ VPWR __dut__._1119_/X sky130_fd_sc_hd__a21o_4
XFILLER_12_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1046__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._0937__A2 prod[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1423_ __dut__.__uuf__._1442_/A VGND VGND VPWR VPWR __dut__.__uuf__._1423_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1354_ __dut__.__uuf__._1380_/A VGND VGND VPWR VPWR __dut__.__uuf__._1354_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1285_ __dut__.__uuf__._1284_/Y __dut__.__uuf__._1276_/X __dut__.__uuf__._1271_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1285_/X sky130_fd_sc_hd__o21a_4
X__dut__._1470_ rst VGND VGND VPWR VPWR __dut__._1470_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0873__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1802__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_280_ _290_/CLK _280_/D VGND VGND VPWR VPWR _280_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_17_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1806_ clkbuf_4_5_0_tck/X __dut__._1806_/D __dut__._1523_/Y VGND VGND VPWR
+ VPWR __dut__._1806_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1737_ __dut__._1543_/Y mp[21] __dut__._1736_/X VGND VGND VPWR VPWR __dut__._1737_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1668_ __dut__._1788_/A __dut__._1821_/Q VGND VGND VPWR VPWR __dut__._1668_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1599_ __dut__._1767_/A1 __dut__._1597_/X __dut__._1598_/X VGND VGND VPWR
+ VPWR __dut__._1803_/D sky130_fd_sc_hd__a21o_4
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1041__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1070_ __dut__.__uuf__._1416_/A VGND VGND VPWR VPWR __dut__.__uuf__._1070_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_67_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1504__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1972_ __dut__._1116_/B VGND VGND VPWR VPWR __dut__.__uuf__._1972_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0970_ __dut__._0970_/A __dut__._1901_/Q VGND VGND VPWR VPWR __dut__._0970_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1406_ __dut__._1218_/B VGND VGND VPWR VPWR __dut__.__uuf__._1406_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1337_ __dut__.__uuf__._1342_/A VGND VGND VPWR VPWR __dut__.__uuf__._1337_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1099__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1522_ rst VGND VGND VPWR VPWR __dut__._1522_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1268_ __dut__.__uuf__._1448_/A VGND VGND VPWR VPWR __dut__.__uuf__._1535_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1453_ rst VGND VGND VPWR VPWR __dut__._1453_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1199_ __dut__.__uuf__._1198_/X __dut__.__uuf__._1195_/X prod[23]
+ prod[24] __dut__.__uuf__._1191_/X VGND VGND VPWR VPWR __dut__._1315_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1384_ __dut__._1542_/A prod[57] VGND VGND VPWR VPWR __dut__._1384_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1414__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ _313_/CLK _263_/D VGND VGND VPWR VPWR _263_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__._1023__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_194_ _194_/A VGND VGND VPWR VPWR _203_/A sky130_fd_sc_hd__inv_2
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1565__A2 mc[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2171_ __dut__.__uuf__._2194_/CLK __dut__._1331_/X __dut__.__uuf__._1172_/X
+ VGND VGND VPWR VPWR prod[31] sky130_fd_sc_hd__dfrtp_4
XFILLER_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1122_ __dut__.__uuf__._1109_/X __dut__.__uuf__._1121_/X prod[49]
+ prod[50] __dut__.__uuf__._1117_/X VGND VGND VPWR VPWR __dut__._1367_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1053_ __dut__._1406_/B __dut__.__uuf__._1057_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1053_/X sky130_fd_sc_hd__or2_4
XFILLER_68_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2109__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1234__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1253__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1955_ __dut__.__uuf__._1951_/Y __dut__.__uuf__._1952_/Y __dut__.__uuf__._1941_/X
+ __dut__.__uuf__._1954_/X VGND VGND VPWR VPWR __dut__.__uuf__._1956_/A sky130_fd_sc_hd__a211o_4
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1886_ __dut__.__uuf__._1941_/A VGND VGND VPWR VPWR __dut__.__uuf__._1886_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._0953_ __dut__._0953_/A1 prod[8] __dut__._0952_/X VGND VGND VPWR VPWR __dut__._1893_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0884_ __dut__._1378_/A __dut__._1858_/Q VGND VGND VPWR VPWR __dut__._0884_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__213__A tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1505_ rst VGND VGND VPWR VPWR __dut__._1505_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_84_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1436_ rst VGND VGND VPWR VPWR __dut__._1436_/Y sky130_fd_sc_hd__inv_2
X__dut__._1367_ __dut__._1383_/A1 __dut__._1367_/A2 __dut__._1366_/X VGND VGND VPWR
+ VPWR __dut__._1367_/X sky130_fd_sc_hd__a21o_4
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1298_ __dut__._1324_/A prod[14] VGND VGND VPWR VPWR __dut__._1298_/X sky130_fd_sc_hd__and2_4
X_315_ _194_/A _315_/D trst VGND VGND VPWR VPWR _315_/Q sky130_fd_sc_hd__dfrtp_4
X_246_ _203_/X _295_/Q VGND VGND VPWR VPWR _246_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_177_ _275_/Q _182_/B VGND VGND VPWR VPWR _274_/D sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_146_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1235__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1740_ __dut__.__uuf__._1773_/A __dut__.__uuf__._1740_/B __dut__.__uuf__._1740_/C
+ VGND VGND VPWR VPWR __dut__._1031_/A2 sky130_fd_sc_hd__and3_4
X__dut__.__uuf__._1671_ __dut__.__uuf__._1573_/X __dut__.__uuf__._1670_/B __dut__.__uuf__._1670_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1672_/C sky130_fd_sc_hd__o21ai_4
Xclkbuf_3_0_0___dut__.__uuf__.__clk_source__ clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_1_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2154_ __dut__.__uuf__._2169_/CLK __dut__._1297_/X __dut__.__uuf__._1222_/X
+ VGND VGND VPWR VPWR prod[14] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1105_ __dut__.__uuf__._1115_/A VGND VGND VPWR VPWR __dut__.__uuf__._1105_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2085_ __dut__.__uuf__._2097_/CLK __dut__._1159_/X __dut__.__uuf__._1529_/X
+ VGND VGND VPWR VPWR __dut__._1160_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_83_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1036_ __dut__.__uuf__._1036_/A __dut__.__uuf__._1036_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1036_/X sky130_fd_sc_hd__or2_4
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1221_ __dut__._1787_/A1 __dut__._1221_/A2 __dut__._1220_/X VGND VGND VPWR
+ VPWR __dut__._1221_/X sky130_fd_sc_hd__a21o_4
X__dut__._1152_ __dut__._1766_/A __dut__._1152_/B VGND VGND VPWR VPWR __dut__._1152_/X
+ sky130_fd_sc_hd__and2_4
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1938_ __dut__.__uuf__._1938_/A __dut__.__uuf__._1938_/B __dut__.__uuf__._1938_/C
+ VGND VGND VPWR VPWR __dut__._1103_/A2 sky130_fd_sc_hd__and3_4
X__dut__._1083_ __dut__._1129_/A1 __dut__._1083_/A2 __dut__._1082_/X VGND VGND VPWR
+ VPWR __dut__._1083_/X sky130_fd_sc_hd__a21o_4
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1777__A2 mp[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1869_ __dut__.__uuf__._1862_/Y __dut__.__uuf__._1863_/Y __dut__.__uuf__._1862_/Y
+ __dut__.__uuf__._1863_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1870_/C sky130_fd_sc_hd__a2bb2o_4
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0936_ __dut__._1404_/A __dut__._0936_/B VGND VGND VPWR VPWR __dut__._0936_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._0867_ __dut__._1767_/A1 __dut__._0865_/X __dut__._0866_/X VGND VGND VPWR
+ VPWR __dut__._1852_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1701__A2 mp[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1419_ rst VGND VGND VPWR VPWR __dut__._1419_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1602__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1217__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_229_ _299_/Q _228_/B _222_/A VGND VGND VPWR VPWR _302_/D sky130_fd_sc_hd__o21a_4
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0888__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1512__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1723_ __dut__.__uuf__._1718_/Y __dut__.__uuf__._1719_/Y __dut__.__uuf__._1686_/X
+ __dut__.__uuf__._1728_/B VGND VGND VPWR VPWR __dut__.__uuf__._1723_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1654_ __dut__.__uuf__._1654_/A VGND VGND VPWR VPWR __dut__.__uuf__._1654_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1585_ __dut__.__uuf__._1587_/A VGND VGND VPWR VPWR __dut__.__uuf__._1585_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1770_ __dut__._1770_/A __dut__._1844_/Q VGND VGND VPWR VPWR __dut__._1770_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._2206_ __dut__.__uuf__._2206_/CLK __dut__._1401_/X __dut__.__uuf__._1060_/X
+ VGND VGND VPWR VPWR __dut__._1402_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1909__CLK __dut__._1917_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2137_ __dut__.__uuf__._2138_/CLK __dut__._1263_/X __dut__.__uuf__._1279_/X
+ VGND VGND VPWR VPWR __dut__._1264_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2068_ __dut__.__uuf__._2119_/CLK __dut__._1125_/X __dut__.__uuf__._1584_/X
+ VGND VGND VPWR VPWR __dut__._1126_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_56_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1019_ __dut__._1400_/B VGND VGND VPWR VPWR __dut__.__uuf__._1029_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_83_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1204_ __dut__._1786_/A __dut__._1204_/B VGND VGND VPWR VPWR __dut__._1204_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1422__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_47_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_104 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1084_/A sky130_fd_sc_hd__buf_2
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_115 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1642_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_126 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1138_/A sky130_fd_sc_hd__buf_2
X__dut__._1135_ __dut__._1787_/A1 __dut__._1135_/A2 __dut__._1134_/X VGND VGND VPWR
+ VPWR __dut__._1135_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_137 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._0940_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_159 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1342_/A sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1054__A __dut__.__uuf__._1100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpsn_inst_psn_buff_148 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1314_/A sky130_fd_sc_hd__buf_2
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1066_ __dut__._1074_/A __dut__._1066_/B VGND VGND VPWR VPWR __dut__._1066_/X
+ sky130_fd_sc_hd__and2_4
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0919_ __dut__._1383_/A1 prod[56] __dut__._0918_/X VGND VGND VPWR VPWR __dut__._1876_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1899_ __dut__._1899_/CLK __dut__._1899_/D __dut__._1430_/Y VGND VGND VPWR
+ VPWR __dut__._1899_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1332__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_109_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__301__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1370_ __dut__.__uuf__._1365_/X __dut__.__uuf__._1369_/X __dut__._1230_/B
+ __dut__.__uuf__._1365_/X VGND VGND VPWR VPWR __dut__._1229_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1677__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1507__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1242__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1601__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1706_ __dut__._1026_/B VGND VGND VPWR VPWR __dut__.__uuf__._1706_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1637_ __dut__.__uuf__._1637_/A VGND VGND VPWR VPWR __dut__.__uuf__._1642_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1822_ clkbuf_4_7_0_tck/X __dut__._1822_/D __dut__._1507_/Y VGND VGND VPWR
+ VPWR __dut__._1822_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1568_ __dut__.__uuf__._1551_/X __dut__.__uuf__._1781_/A __dut__._1142_/B
+ __dut__.__uuf__._1449_/A __dut__.__uuf__._1567_/X VGND VGND VPWR VPWR __dut__._1141_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1499_ __dut__._1717_/X __dut__.__uuf__._1494_/X __dut__._1178_/B
+ __dut__.__uuf__._1495_/X VGND VGND VPWR VPWR __dut__.__uuf__._1499_/X sky130_fd_sc_hd__o22a_4
X__dut__._1753_ __dut__._1543_/Y mp[25] __dut__._1752_/X VGND VGND VPWR VPWR __dut__._1753_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1684_ __dut__._1788_/A __dut__._1825_/Q VGND VGND VPWR VPWR __dut__._1684_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_88_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1417__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1152__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1118_ __dut__._1678_/A __dut__._1118_/B VGND VGND VPWR VPWR __dut__._1118_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1049_ __dut__._1049_/A1 __dut__._1049_/A2 __dut__._1048_/X VGND VGND VPWR
+ VPWR __dut__._1049_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1659__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1062__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__.__uuf__._2142__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1422_ __dut__.__uuf__._1469_/A VGND VGND VPWR VPWR __dut__.__uuf__._1442_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1353_ __dut__.__uuf__._1367_/A VGND VGND VPWR VPWR __dut__.__uuf__._1353_/X
+ sky130_fd_sc_hd__buf_2
Xclkbuf_4_3_0_tck clkbuf_4_3_0_tck/A VGND VGND VPWR VPWR _194_/A sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1284_ __dut__._1264_/B VGND VGND VPWR VPWR __dut__.__uuf__._1284_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._0873__A2 mc[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__294__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1700__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1805_ clkbuf_4_5_0_tck/X __dut__._1805_/D __dut__._1524_/Y VGND VGND VPWR
+ VPWR __dut__._1805_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._2015__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1736_ __dut__._1788_/A __dut__._1838_/Q VGND VGND VPWR VPWR __dut__._1736_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_1_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1667_ __dut__._1767_/A1 __dut__._1665_/X __dut__._1666_/X VGND VGND VPWR
+ VPWR __dut__._1820_/D sky130_fd_sc_hd__a21o_4
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0986__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1598_ __dut__._1766_/A __dut__._1802_/Q VGND VGND VPWR VPWR __dut__._1598_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1610__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0896__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1971_ __dut__._1122_/B VGND VGND VPWR VPWR __dut__.__uuf__._1971_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_23_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1520__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2038__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1405_ __dut__.__uuf__._1416_/A VGND VGND VPWR VPWR __dut__.__uuf__._1405_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1336_ __dut__.__uuf__._1329_/X __dut__.__uuf__._1335_/X __dut__._1244_/B
+ __dut__.__uuf__._1329_/X VGND VGND VPWR VPWR __dut__._1243_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1521_ rst VGND VGND VPWR VPWR __dut__._1521_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1267_ __dut__._1268_/B VGND VGND VPWR VPWR __dut__.__uuf__._1267_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1452_ rst VGND VGND VPWR VPWR __dut__._1452_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1198_ __dut__.__uuf__._1212_/A VGND VGND VPWR VPWR __dut__.__uuf__._1198_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1383_ __dut__._1383_/A1 __dut__._1383_/A2 __dut__._1382_/X VGND VGND VPWR
+ VPWR __dut__._1383_/X sky130_fd_sc_hd__a21o_4
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1430__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_262_ _314_/CLK _262_/D VGND VGND VPWR VPWR _262_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA___dut__.__uuf__._1091__B1 prod[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_193_ _260_/Q _193_/B VGND VGND VPWR VPWR _259_/D sky130_fd_sc_hd__or2_4
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1719_ __dut__._1719_/A1 __dut__._1717_/X __dut__._1718_/X VGND VGND VPWR
+ VPWR __dut__._1833_/D sky130_fd_sc_hd__a21o_4
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2170_ __dut__.__uuf__._2194_/CLK __dut__._1329_/X __dut__.__uuf__._1174_/X
+ VGND VGND VPWR VPWR prod[30] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1121_ __dut__.__uuf__._1149_/A VGND VGND VPWR VPWR __dut__.__uuf__._1121_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_87_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1052_ __dut__.__uuf__._1052_/A VGND VGND VPWR VPWR __dut__.__uuf__._1052_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1515__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1954_ __dut__.__uuf__._1951_/Y __dut__.__uuf__._1952_/Y __dut__.__uuf__._1908_/X
+ __dut__.__uuf__._1958_/B VGND VGND VPWR VPWR __dut__.__uuf__._1954_/X sky130_fd_sc_hd__o22a_4
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1885_ __dut__._1084_/B VGND VGND VPWR VPWR __dut__.__uuf__._1885_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._0952_ __dut__._1770_/A __dut__._1892_/Q VGND VGND VPWR VPWR __dut__._0952_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0883_ __dut__._0883_/A1 prod[38] __dut__._0882_/X VGND VGND VPWR VPWR __dut__._1858_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_87_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1319_ __dut__.__uuf__._1314_/X __dut__.__uuf__._1318_/X __dut__._1250_/B
+ __dut__.__uuf__._1314_/X VGND VGND VPWR VPWR __dut__._1249_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__._1504_ rst VGND VGND VPWR VPWR __dut__._1504_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1425__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_77_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1435_ rst VGND VGND VPWR VPWR __dut__._1435_/Y sky130_fd_sc_hd__inv_2
X__dut__._1366_ __dut__._1378_/A prod[48] VGND VGND VPWR VPWR __dut__._1366_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2203__CLK __dut__.__uuf__._2210_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1297_ __dut__._1319_/A1 __dut__._1297_/A2 __dut__._1296_/X VGND VGND VPWR
+ VPWR __dut__._1297_/X sky130_fd_sc_hd__a21o_4
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1160__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_314_ _314_/CLK _314_/D trst VGND VGND VPWR VPWR _314_/Q sky130_fd_sc_hd__dfrtp_4
X_245_ tdi _154_/C _302_/Q _315_/Q VGND VGND VPWR VPWR _315_/D sky130_fd_sc_hd__o22a_4
XFILLER_6_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_176_ _183_/A VGND VGND VPWR VPWR _182_/B sky130_fd_sc_hd__buf_2
XFILLER_69_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_139_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1670_ __dut__.__uuf__._1692_/A __dut__.__uuf__._1670_/B __dut__.__uuf__._1670_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1672_/B sky130_fd_sc_hd__or3_4
XANTENNA___dut__._1171__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2153_ __dut__.__uuf__._2169_/CLK __dut__._1295_/X __dut__.__uuf__._1225_/X
+ VGND VGND VPWR VPWR prod[13] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1104_ __dut__.__uuf__._1162_/A VGND VGND VPWR VPWR __dut__.__uuf__._1115_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_87_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2084_ __dut__.__uuf__._2097_/CLK __dut__._1157_/X __dut__.__uuf__._1534_/X
+ VGND VGND VPWR VPWR __dut__._1158_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_83_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1035_ __dut__.__uuf__._1037_/B VGND VGND VPWR VPWR __dut__.__uuf__._1036_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._1220_ __dut__._1786_/A __dut__._1220_/B VGND VGND VPWR VPWR __dut__._1220_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1151_ __dut__._1151_/A1 __dut__._1151_/A2 __dut__._1150_/X VGND VGND VPWR
+ VPWR __dut__._1151_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1937_ __dut__.__uuf__._1936_/X __dut__.__uuf__._1935_/B __dut__.__uuf__._1935_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1938_/C sky130_fd_sc_hd__o21ai_4
X__dut__._1082_ __dut__._1082_/A __dut__._1082_/B VGND VGND VPWR VPWR __dut__._1082_/X
+ sky130_fd_sc_hd__and2_4
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1868_ __dut__.__uuf__._1868_/A VGND VGND VPWR VPWR __dut__.__uuf__._1914_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1838__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1799_ __dut__._1581_/X VGND VGND VPWR VPWR __dut__.__uuf__._1804_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._0935_ __dut__._1405_/A1 done __dut__._0934_/X VGND VGND VPWR VPWR __dut__._1884_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0866_ __dut__._1766_/A __dut__._1851_/Q VGND VGND VPWR VPWR __dut__._0866_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0994__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1418_ rst VGND VGND VPWR VPWR __dut__._1418_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1349_ __dut__._1349_/A1 __dut__._1349_/A2 __dut__._1348_/X VGND VGND VPWR
+ VPWR __dut__._1349_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._1515__A __dut__.__uuf__._1536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_228_ _232_/A _228_/B VGND VGND VPWR VPWR _301_/D sky130_fd_sc_hd__and2_4
X_159_ _289_/Q _164_/B VGND VGND VPWR VPWR _288_/D sky130_fd_sc_hd__and2_4
XFILLER_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1722_ __dut__._1613_/X VGND VGND VPWR VPWR __dut__.__uuf__._1728_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1653_ __dut__.__uuf__._1654_/A VGND VGND VPWR VPWR __dut__.__uuf__._1653_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1584_ __dut__.__uuf__._1587_/A VGND VGND VPWR VPWR __dut__.__uuf__._1584_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2205_ __dut__.__uuf__._2210_/CLK __dut__._1399_/X __dut__.__uuf__._1063_/X
+ VGND VGND VPWR VPWR __dut__._1400_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_0_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._2136_ __dut__.__uuf__._2138_/CLK __dut__._1261_/X __dut__.__uuf__._1283_/X
+ VGND VGND VPWR VPWR __dut__._1262_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2067_ __dut__.__uuf__._2119_/CLK __dut__._1123_/X __dut__.__uuf__._1585_/X
+ VGND VGND VPWR VPWR __dut__._1124_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1018_ __dut__._1136_/B VGND VGND VPWR VPWR __dut__.__uuf__._2005_/A
+ sky130_fd_sc_hd__inv_2
XFILLER_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1203_ __dut__._1779_/A1 __dut__._1203_/A2 __dut__._1202_/X VGND VGND VPWR
+ VPWR __dut__._1203_/X sky130_fd_sc_hd__a21o_4
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_105 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1082_/A sky130_fd_sc_hd__buf_2
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_116 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1146_/A sky130_fd_sc_hd__buf_2
X__dut__._1134_ __dut__._1786_/A __dut__._1134_/B VGND VGND VPWR VPWR __dut__._1134_/X
+ sky130_fd_sc_hd__and2_4
Xpsn_inst_psn_buff_127 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1180_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_149 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1316_/A sky130_fd_sc_hd__buf_2
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1065_ __dut__._1071_/A1 __dut__._1065_/A2 __dut__._1064_/X VGND VGND VPWR
+ VPWR __dut__._1065_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_138 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._0942_/A sky130_fd_sc_hd__buf_2
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1383__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0918_ __dut__._1542_/A __dut__._1875_/Q VGND VGND VPWR VPWR __dut__._0918_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1135__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1898_ __dut__._1899_/CLK __dut__._1898_/D __dut__._1431_/Y VGND VGND VPWR
+ VPWR __dut__._1898_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._2071__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1677__A2 mc[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1523__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1264__A3 prod[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1601__A2 mc[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1705_ __dut__.__uuf__._1717_/A __dut__.__uuf__._1705_/B __dut__.__uuf__._1705_/C
+ VGND VGND VPWR VPWR __dut__._1019_/A2 sky130_fd_sc_hd__and3_4
X__dut__.__uuf__._1636_ __dut__.__uuf__._1636_/A VGND VGND VPWR VPWR __dut__.__uuf__._1636_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1365__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1821_ clkbuf_4_7_0_tck/X __dut__._1821_/D __dut__._1508_/Y VGND VGND VPWR
+ VPWR __dut__._1821_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1567_ __dut__._1645_/X __dut__.__uuf__._1078_/A __dut__._1144_/B
+ __dut__.__uuf__._1660_/A VGND VGND VPWR VPWR __dut__.__uuf__._1567_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__._1117__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1498_ __dut__.__uuf__._1508_/A VGND VGND VPWR VPWR __dut__.__uuf__._1498_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1752_ __dut__._1788_/A __dut__._1842_/Q VGND VGND VPWR VPWR __dut__._1752_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1683_ __dut__._1767_/A1 __dut__._1681_/X __dut__._1682_/X VGND VGND VPWR
+ VPWR __dut__._1824_/D sky130_fd_sc_hd__a21o_4
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2119_ __dut__.__uuf__._2119_/CLK __dut__._1227_/X __dut__.__uuf__._1373_/X
+ VGND VGND VPWR VPWR __dut__._1228_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_29_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1433__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1117_ __dut__._1129_/A1 __dut__._1117_/A2 __dut__._1116_/X VGND VGND VPWR
+ VPWR __dut__._1117_/X sky130_fd_sc_hd__a21o_4
XFILLER_8_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1048_ __dut__._1678_/A __dut__._1048_/B VGND VGND VPWR VPWR __dut__._1048_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__.__uuf__._2094__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1608__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_121_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1595__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1421_ __dut__.__uuf__._1416_/X __dut__.__uuf__._1420_/X __dut__._1210_/B
+ __dut__.__uuf__._1416_/X VGND VGND VPWR VPWR __dut__._1209_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1352_ __dut__.__uuf__._1340_/X __dut__.__uuf__._1351_/X __dut__._1238_/B
+ __dut__.__uuf__._1340_/X VGND VGND VPWR VPWR __dut__._1237_/A2 sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._1518__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1283_ __dut__.__uuf__._1288_/A VGND VGND VPWR VPWR __dut__.__uuf__._1283_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1619_ __dut__.__uuf__._1637_/A VGND VGND VPWR VPWR __dut__.__uuf__._1624_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1804_ clkbuf_4_5_0_tck/X __dut__._1804_/D __dut__._1525_/Y VGND VGND VPWR
+ VPWR __dut__._1804_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1735_ __dut__._1735_/A1 __dut__._1733_/X __dut__._1734_/X VGND VGND VPWR
+ VPWR __dut__._1837_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1428__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1666_ __dut__._1766_/A __dut__._1819_/Q VGND VGND VPWR VPWR __dut__._1666_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1597_ __dut__._1543_/Y mc[21] __dut__._1596_/X VGND VGND VPWR VPWR __dut__._1597_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1577__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_169_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1970_ __dut__.__uuf__._1990_/A __dut__.__uuf__._1970_/B __dut__.__uuf__._1970_/C
+ VGND VGND VPWR VPWR __dut__._1115_/A2 sky130_fd_sc_hd__and3_4
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1871__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1404_ __dut__.__uuf__._1418_/A VGND VGND VPWR VPWR __dut__.__uuf__._1404_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1335_ __dut__.__uuf__._1334_/Y __dut__.__uuf__._1323_/X __dut__.__uuf__._1324_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1335_/X sky130_fd_sc_hd__o21a_4
X__dut__._1520_ rst VGND VGND VPWR VPWR __dut__._1520_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1266_ __dut__.__uuf__._1288_/A VGND VGND VPWR VPWR __dut__.__uuf__._1266_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1451_ rst VGND VGND VPWR VPWR __dut__._1451_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1197_ __dut__.__uuf__._1204_/A VGND VGND VPWR VPWR __dut__.__uuf__._1197_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1382_ __dut__._1542_/A prod[56] VGND VGND VPWR VPWR __dut__._1382_/X sky130_fd_sc_hd__and2_4
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1559__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_261_ _313_/CLK _261_/D VGND VGND VPWR VPWR _261_/Q sky130_fd_sc_hd__dfxtp_4
X_192_ _261_/Q _193_/B VGND VGND VPWR VPWR _260_/D sky130_fd_sc_hd__or2_4
XANTENNA_psn_inst_psn_buff_22_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1158__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1718_ __dut__._1766_/A __dut__._1832_/Q VGND VGND VPWR VPWR __dut__._1718_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1649_ __dut__._1543_/Y mp[1] __dut__._1648_/X VGND VGND VPWR VPWR __dut__._1649_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_2_0_tck clkbuf_4_3_0_tck/A VGND VGND VPWR VPWR _314_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_60_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1894__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1120_ __dut__.__uuf__._1130_/A VGND VGND VPWR VPWR __dut__.__uuf__._1120_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_87_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1051_ __dut__.__uuf__._1063_/A VGND VGND VPWR VPWR __dut__.__uuf__._1051_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_83_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1789__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1953_ __dut__._1721_/X VGND VGND VPWR VPWR __dut__.__uuf__._1958_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_24_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1531__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1884_ __dut__._1090_/B VGND VGND VPWR VPWR __dut__.__uuf__._1884_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._0951_ __dut__._0951_/A1 prod[7] __dut__._0950_/X VGND VGND VPWR VPWR __dut__._1892_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0882_ __dut__._0882_/A __dut__._1857_/Q VGND VGND VPWR VPWR __dut__._0882_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1713__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1318_ __dut__.__uuf__._1317_/Y __dut__.__uuf__._1297_/X __dut__.__uuf__._1299_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1318_/X sky130_fd_sc_hd__o21a_4
X__dut__._1503_ rst VGND VGND VPWR VPWR __dut__._1503_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1706__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1249_ __dut__.__uuf__._1249_/A VGND VGND VPWR VPWR __dut__.__uuf__._1249_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_59_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1434_ rst VGND VGND VPWR VPWR __dut__._1434_/Y sky130_fd_sc_hd__inv_2
X__dut__._1365_ __dut__._1383_/A1 __dut__._1365_/A2 __dut__._1364_/X VGND VGND VPWR
+ VPWR __dut__._1365_/X sky130_fd_sc_hd__a21o_4
X__dut__._1296_ __dut__._1770_/A prod[13] VGND VGND VPWR VPWR __dut__._1296_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1441__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_313_ _313_/CLK _313_/D trst VGND VGND VPWR VPWR _313_/Q sky130_fd_sc_hd__dfrtp_4
X_244_ _312_/Q _311_/Q _244_/C _244_/D VGND VGND VPWR VPWR _244_/X sky130_fd_sc_hd__and4_4
XFILLER_6_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_175_ _276_/Q _187_/B VGND VGND VPWR VPWR _275_/D sky130_fd_sc_hd__or2_4
XANTENNA___dut__._1616__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2028__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__309__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2152_ __dut__.__uuf__._2169_/CLK __dut__._1293_/X __dut__.__uuf__._1229_/X
+ VGND VGND VPWR VPWR prod[12] sky130_fd_sc_hd__dfrtp_4
XFILLER_87_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1103_ __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR __dut__.__uuf__._1162_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1526__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2083_ __dut__.__uuf__._2083_/CLK __dut__._1155_/X __dut__.__uuf__._1540_/X
+ VGND VGND VPWR VPWR __dut__._1156_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1034_ __dut__._1408_/B __dut__.__uuf__._1052_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1037_/B sky130_fd_sc_hd__and2_4
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1150_ __dut__._1150_/A __dut__._1150_/B VGND VGND VPWR VPWR __dut__._1150_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_36_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1936_ __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR __dut__.__uuf__._1936_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1081_ __dut__._1129_/A1 __dut__._1081_/A2 __dut__._1080_/X VGND VGND VPWR
+ VPWR __dut__._1081_/X sky130_fd_sc_hd__a21o_4
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1867_ __dut__.__uuf__._1867_/A VGND VGND VPWR VPWR __dut__._1081_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1798_ __dut__.__uuf__._1923_/A VGND VGND VPWR VPWR __dut__.__uuf__._1798_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0934_ __dut__._1408_/A __dut__._1883_/Q VGND VGND VPWR VPWR __dut__._0934_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._0865_ __dut__._1543_/Y mc[7] __dut__._0864_/X VGND VGND VPWR VPWR __dut__._0865_/X
+ sky130_fd_sc_hd__a21o_4
Xclkbuf_2_2_0___dut__.__uuf__.__clk_source__ clkbuf_2_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1436__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1417_ rst VGND VGND VPWR VPWR __dut__._1417_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1348_ __dut__._1378_/A prod[39] VGND VGND VPWR VPWR __dut__._1348_/X sky130_fd_sc_hd__and2_4
XFILLER_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1279_ __dut__._1279_/A1 __dut__._1279_/A2 __dut__._1278_/X VGND VGND VPWR
+ VPWR __dut__._1279_/X sky130_fd_sc_hd__a21o_4
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_227_ _302_/Q _303_/Q VGND VGND VPWR VPWR _228_/B sky130_fd_sc_hd__or2_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_158_ _290_/Q _164_/B VGND VGND VPWR VPWR _289_/D sky130_fd_sc_hd__and2_4
XFILLER_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_151_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1721_ __dut__.__uuf__._1941_/A VGND VGND VPWR VPWR __dut__.__uuf__._1721_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1652_ __dut__.__uuf__._1654_/A VGND VGND VPWR VPWR __dut__.__uuf__._1652_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA__281__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1583_ __dut__.__uuf__._1587_/A VGND VGND VPWR VPWR __dut__.__uuf__._1583_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2204_ __dut__.__uuf__._2210_/CLK __dut__._1397_/X __dut__.__uuf__._1068_/X
+ VGND VGND VPWR VPWR __dut__._1398_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1256__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2135_ __dut__.__uuf__._2138_/CLK __dut__._1259_/X __dut__.__uuf__._1288_/X
+ VGND VGND VPWR VPWR __dut__._1260_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2066_ __dut__.__uuf__._2119_/CLK __dut__._1121_/X __dut__.__uuf__._1586_/X
+ VGND VGND VPWR VPWR __dut__._1122_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1805__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1202_ __dut__._1786_/A __dut__._1202_/B VGND VGND VPWR VPWR __dut__._1202_/X
+ sky130_fd_sc_hd__and2_4
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_106 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1054_/A sky130_fd_sc_hd__buf_2
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_117 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1144_/A sky130_fd_sc_hd__buf_2
X__dut__._1133_ __dut__._1787_/A1 __dut__._1133_/A2 __dut__._1132_/X VGND VGND VPWR
+ VPWR __dut__._1133_/X sky130_fd_sc_hd__a21o_4
Xpsn_inst_psn_buff_128 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1188_/A sky130_fd_sc_hd__buf_2
XFILLER_12_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1919_ __dut__._0865_/X VGND VGND VPWR VPWR __dut__.__uuf__._1925_/B
+ sky130_fd_sc_hd__inv_2
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1064_ __dut__._1074_/A __dut__._1064_/B VGND VGND VPWR VPWR __dut__._1064_/X
+ sky130_fd_sc_hd__and2_4
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_139 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._0974_/A sky130_fd_sc_hd__buf_2
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__235__A _251_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0917_ __dut__._1383_/A1 prod[55] __dut__._0916_/X VGND VGND VPWR VPWR __dut__._1875_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1897_ __dut__._1899_/CLK __dut__._1897_/D __dut__._1432_/Y VGND VGND VPWR
+ VPWR __dut__._1897_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1166__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1076__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__310__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1704_ __dut__.__uuf__._1573_/X __dut__.__uuf__._1703_/B __dut__.__uuf__._1703_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1705_/C sky130_fd_sc_hd__o21ai_4
X__dut__.__uuf__._1635_ __dut__.__uuf__._1636_/A VGND VGND VPWR VPWR __dut__.__uuf__._1635_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1820_ clkbuf_4_7_0_tck/X __dut__._1820_/D __dut__._1509_/Y VGND VGND VPWR
+ VPWR __dut__._1820_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1566_ __dut__.__uuf__._1566_/A VGND VGND VPWR VPWR __dut__.__uuf__._1781_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1497_ __dut__.__uuf__._1487_/X __dut__.__uuf__._1483_/X __dut__._1178_/B
+ __dut__.__uuf__._1493_/X __dut__.__uuf__._1496_/X VGND VGND VPWR VPWR __dut__._1177_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1751_ __dut__._1759_/A1 __dut__._1749_/X __dut__._1750_/X VGND VGND VPWR
+ VPWR __dut__._1841_/D sky130_fd_sc_hd__a21o_4
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1682_ __dut__._1766_/A __dut__._1822_/Q VGND VGND VPWR VPWR __dut__._1682_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2118_ __dut__.__uuf__._2119_/CLK __dut__._1225_/X __dut__.__uuf__._1379_/X
+ VGND VGND VPWR VPWR __dut__._1226_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2049_ __dut__.__uuf__._2049_/CLK __dut__._1087_/X __dut__.__uuf__._1607_/X
+ VGND VGND VPWR VPWR __dut__._1088_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1714__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_52_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1116_ __dut__._1116_/A __dut__._1116_/B VGND VGND VPWR VPWR __dut__._1116_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1047_ __dut__._1047_/A1 __dut__._1047_/A2 __dut__._1046_/X VGND VGND VPWR
+ VPWR __dut__._1047_/X sky130_fd_sc_hd__a21o_4
XFILLER_40_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0867__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1624__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_114_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__145__A3 tdi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1420_ __dut__.__uuf__._1419_/Y __dut__.__uuf__._1400_/X __dut__.__uuf__._1401_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1420_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1351_ __dut__.__uuf__._1348_/Y __dut__.__uuf__._1349_/X __dut__.__uuf__._1350_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1351_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1282_ __dut__.__uuf__._1274_/X __dut__.__uuf__._1281_/X __dut__._1264_/B
+ __dut__.__uuf__._1274_/X VGND VGND VPWR VPWR __dut__._1263_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1534__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1035__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1618_ __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR __dut__.__uuf__._1618_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1803_ clkbuf_4_5_0_tck/X __dut__._1803_/D __dut__._1526_/Y VGND VGND VPWR
+ VPWR __dut__._1803_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1549_ __dut__.__uuf__._1530_/X __dut__.__uuf__._1547_/X __dut__._1152_/B
+ __dut__.__uuf__._1535_/X __dut__.__uuf__._1548_/X VGND VGND VPWR VPWR __dut__._1151_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_89_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1734_ __dut__._1770_/A __dut__._1836_/Q VGND VGND VPWR VPWR __dut__._1734_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1665_ __dut__._1543_/Y mp[5] __dut__._1664_/X VGND VGND VPWR VPWR __dut__._1665_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1596_ __dut__._1788_/A __dut__._1803_/Q VGND VGND VPWR VPWR __dut__._1596_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1444__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1577__A2 mc[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1354__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1265__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1017__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1529__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1403_ __dut__.__uuf__._1391_/X __dut__.__uuf__._1402_/X __dut__._1218_/B
+ __dut__.__uuf__._1391_/X VGND VGND VPWR VPWR __dut__._1217_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1334_ __dut__._1246_/B VGND VGND VPWR VPWR __dut__.__uuf__._1334_/Y
+ sky130_fd_sc_hd__inv_2
Xclkbuf_4_3_0___dut__.__uuf__.__clk_source__ clkbuf_4_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2114_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1265_ __dut__.__uuf__._1346_/A VGND VGND VPWR VPWR __dut__.__uuf__._1288_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_58_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1450_ rst VGND VGND VPWR VPWR __dut__._1450_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1196_ __dut__.__uuf__._1183_/X __dut__.__uuf__._1195_/X prod[24]
+ prod[25] __dut__.__uuf__._1191_/X VGND VGND VPWR VPWR __dut__._1317_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1381_ __dut__._1383_/A1 __dut__._1381_/A2 __dut__._1380_/X VGND VGND VPWR
+ VPWR __dut__._1381_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1264__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1559__A2 __dut__._1557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_260_ _194_/A _260_/D VGND VGND VPWR VPWR _260_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_191_ _262_/Q _191_/B VGND VGND VPWR VPWR _261_/D sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_15_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1439__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1717_ __dut__._1543_/Y mp[17] __dut__._1716_/X VGND VGND VPWR VPWR __dut__._1717_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1648_ __dut__._1788_/A __dut__._1816_/Q VGND VGND VPWR VPWR __dut__._1648_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1579_ __dut__._1767_/A1 __dut__._1577_/X __dut__._1578_/X VGND VGND VPWR
+ VPWR __dut__._1798_/D sky130_fd_sc_hd__a21o_4
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1247__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1050_ __dut__.__uuf__._1100_/A __dut__.__uuf__._1049_/X __dut__.__uuf__._1036_/B
+ __dut__._1408_/B __dut__.__uuf__._1043_/X VGND VGND VPWR VPWR __dut__._1407_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_68_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1789__A2 mc[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1952_ __dut__._1108_/B VGND VGND VPWR VPWR __dut__.__uuf__._1952_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1883_ __dut__.__uuf__._1883_/A __dut__.__uuf__._1883_/B __dut__.__uuf__._1883_/C
+ VGND VGND VPWR VPWR __dut__._1083_/A2 sky130_fd_sc_hd__and3_4
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._0950_ __dut__._1770_/A __dut__._1891_/Q VGND VGND VPWR VPWR __dut__._0950_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._0881_ __dut__._0881_/A1 prod[37] __dut__._0880_/X VGND VGND VPWR VPWR __dut__._1857_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1713__A2 mp[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1317_ __dut__._1252_/B VGND VGND VPWR VPWR __dut__.__uuf__._1317_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_59_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1502_ rst VGND VGND VPWR VPWR __dut__._1502_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1248_ __dut__.__uuf__._1248_/A VGND VGND VPWR VPWR __dut__.__uuf__._1248_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1179_ __dut__.__uuf__._1189_/A VGND VGND VPWR VPWR __dut__.__uuf__._1179_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1433_ rst VGND VGND VPWR VPWR __dut__._1433_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1364_ __dut__._1378_/A prod[47] VGND VGND VPWR VPWR __dut__._1364_/X sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1722__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1229__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1295_ __dut__._1295_/A1 __dut__._1295_/A2 __dut__._1294_/X VGND VGND VPWR
+ VPWR __dut__._1295_/X sky130_fd_sc_hd__a21o_4
X_312_ _194_/A _312_/D trst VGND VGND VPWR VPWR _312_/Q sky130_fd_sc_hd__dfstp_4
X_243_ _301_/Q _300_/Q _302_/Q VGND VGND VPWR VPWR _244_/D sky130_fd_sc_hd__or3_4
XANTENNA___dut__._1401__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_174_ _193_/B VGND VGND VPWR VPWR _187_/B sky130_fd_sc_hd__buf_2
XFILLER_96_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1861__CLK __dut__._1917_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1632__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2151_ __dut__.__uuf__._2169_/CLK __dut__._1291_/X __dut__.__uuf__._1231_/X
+ VGND VGND VPWR VPWR prod[11] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2082_ __dut__.__uuf__._2097_/CLK __dut__._1153_/X __dut__.__uuf__._1543_/X
+ VGND VGND VPWR VPWR __dut__._1154_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1102_ __dut__.__uuf__._1102_/A VGND VGND VPWR VPWR __dut__.__uuf__._1649_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1439__A __dut__.__uuf__._1536_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1033_ __dut__._1406_/B __dut__.__uuf__._1057_/A VGND VGND VPWR VPWR
+ __dut__.__uuf__._1052_/A sky130_fd_sc_hd__and2_4
XFILLER_95_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1542__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1935_ __dut__.__uuf__._1968_/A __dut__.__uuf__._1935_/B __dut__.__uuf__._1935_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1938_/B sky130_fd_sc_hd__or3_4
X__dut__._1080_ __dut__._1678_/A __dut__._1080_/B VGND VGND VPWR VPWR __dut__._1080_/X
+ sky130_fd_sc_hd__and2_4
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1631__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1866_ __dut__.__uuf__._1862_/Y __dut__.__uuf__._1863_/Y __dut__.__uuf__._1831_/X
+ __dut__.__uuf__._1865_/X VGND VGND VPWR VPWR __dut__.__uuf__._1867_/A sky130_fd_sc_hd__a211o_4
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1797_ __dut__._1052_/B VGND VGND VPWR VPWR __dut__.__uuf__._1797_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._0933_ __dut__._1409_/A1 prod[63] __dut__._0932_/X VGND VGND VPWR VPWR __dut__._1883_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0864_ __dut__._1788_/A __dut__._1852_/Q VGND VGND VPWR VPWR __dut__._0864_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_1_0_tck clkbuf_4_1_0_tck/A VGND VGND VPWR VPWR _306_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1884__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_82_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1416_ rst VGND VGND VPWR VPWR __dut__._1416_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1452__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1347_ __dut__._1349_/A1 __dut__._1347_/A2 __dut__._1346_/X VGND VGND VPWR
+ VPWR __dut__._1347_/X sky130_fd_sc_hd__a21o_4
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1278_ __dut__._1280_/A prod[4] VGND VGND VPWR VPWR __dut__._1278_/X sky130_fd_sc_hd__and2_4
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_226_ _301_/Q _300_/Q _222_/A VGND VGND VPWR VPWR _300_/D sky130_fd_sc_hd__o21a_4
X_157_ tdi _164_/B VGND VGND VPWR VPWR _290_/D sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1689__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_144_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1362__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2145__CLK __dut__.__uuf__._2164_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1613__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1720_ __dut__.__uuf__._1720_/A VGND VGND VPWR VPWR __dut__.__uuf__._1941_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1651_ __dut__.__uuf__._1654_/A VGND VGND VPWR VPWR __dut__.__uuf__._1651_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1582_ __dut__.__uuf__._1606_/A VGND VGND VPWR VPWR __dut__.__uuf__._1587_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2203_ __dut__.__uuf__._2210_/CLK __dut__._1395_/X __dut__.__uuf__._1072_/X
+ VGND VGND VPWR VPWR prod[63] sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1537__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2134_ __dut__.__uuf__._2138_/CLK __dut__._1257_/X __dut__.__uuf__._1293_/X
+ VGND VGND VPWR VPWR __dut__._1258_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2065_ __dut__.__uuf__._2065_/CLK __dut__._1119_/X __dut__.__uuf__._1587_/X
+ VGND VGND VPWR VPWR __dut__._1120_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1201_ __dut__._1779_/A1 __dut__._1201_/A2 __dut__._1200_/X VGND VGND VPWR
+ VPWR __dut__._1201_/X sky130_fd_sc_hd__a21o_4
XFILLER_83_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpsn_inst_psn_buff_107 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1056_/A sky130_fd_sc_hd__buf_2
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xpsn_inst_psn_buff_118 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1142_/A sky130_fd_sc_hd__buf_2
X__dut__._1132_ __dut__._1786_/A __dut__._1132_/B VGND VGND VPWR VPWR __dut__._1132_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1918_ __dut__._1096_/B VGND VGND VPWR VPWR __dut__.__uuf__._1918_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1063_ __dut__._1767_/A1 __dut__._1063_/A2 __dut__._1062_/X VGND VGND VPWR
+ VPWR __dut__._1063_/X sky130_fd_sc_hd__a21o_4
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_129 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1190_/A sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1849_ __dut__.__uuf__._1826_/X __dut__.__uuf__._1848_/B __dut__.__uuf__._1848_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1850_/C sky130_fd_sc_hd__o21ai_4
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._0916_ __dut__._1542_/A __dut__._1874_/Q VGND VGND VPWR VPWR __dut__._0916_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2018__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1447__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1896_ __dut__._1899_/CLK __dut__._1896_/D __dut__._1433_/Y VGND VGND VPWR
+ VPWR __dut__._1896_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1182__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_209_ _247_/Q VGND VGND VPWR VPWR _209_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1703_ __dut__.__uuf__._1749_/A __dut__.__uuf__._1703_/B __dut__.__uuf__._1703_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1705_/B sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1634_ __dut__.__uuf__._1636_/A VGND VGND VPWR VPWR __dut__.__uuf__._1634_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1565_ __dut__.__uuf__._1569_/A VGND VGND VPWR VPWR __dut__.__uuf__._1565_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1750_ __dut__._1770_/A __dut__._1840_/Q VGND VGND VPWR VPWR __dut__._1750_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1496_ __dut__._1725_/X __dut__.__uuf__._1494_/X __dut__._1180_/B
+ __dut__.__uuf__._1495_/X VGND VGND VPWR VPWR __dut__.__uuf__._1496_/X sky130_fd_sc_hd__o22a_4
X__dut__._1681_ __dut__._1543_/Y mp[8] __dut__._1680_/X VGND VGND VPWR VPWR __dut__._1681_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_95_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2117_ __dut__.__uuf__._2119_/CLK __dut__._1223_/X __dut__.__uuf__._1384_/X
+ VGND VGND VPWR VPWR __dut__._1224_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2048_ __dut__.__uuf__._2049_/CLK __dut__._1085_/X __dut__.__uuf__._1608_/X
+ VGND VGND VPWR VPWR __dut__._1086_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_45_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1115_ __dut__._1129_/A1 __dut__._1115_/A2 __dut__._1114_/X VGND VGND VPWR
+ VPWR __dut__._1115_/X sky130_fd_sc_hd__a21o_4
XFILLER_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1730__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1046_ __dut__._1678_/A __dut__._1046_/B VGND VGND VPWR VPWR __dut__._1046_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1879_ __dut__._1919_/CLK __dut__._1879_/D __dut__._1450_/Y VGND VGND VPWR
+ VPWR __dut__._1879_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._0867__A2 __dut__._0865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1537__A __dut__.__uuf__._1720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__271__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1640__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_107_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1350_ __dut__.__uuf__._1401_/A VGND VGND VPWR VPWR __dut__.__uuf__._1350_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1281_ __dut__.__uuf__._1280_/Y __dut__.__uuf__._1276_/X __dut__.__uuf__._1271_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1281_/X sky130_fd_sc_hd__o21a_4
XFILLER_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1550__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1617_ __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR __dut__.__uuf__._1617_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1802_ clkbuf_4_5_0_tck/X __dut__._1802_/D __dut__._1527_/Y VGND VGND VPWR
+ VPWR __dut__._1802_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1548_ __dut__._1665_/X __dut__.__uuf__._1536_/X __dut__._1154_/B
+ __dut__.__uuf__._1537_/X VGND VGND VPWR VPWR __dut__.__uuf__._1548_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1479_ __dut__.__uuf__._1486_/A VGND VGND VPWR VPWR __dut__.__uuf__._1479_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1733_ __dut__._1543_/Y mp[20] __dut__._1732_/X VGND VGND VPWR VPWR __dut__._1733_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1664_ __dut__._1788_/A __dut__._1820_/Q VGND VGND VPWR VPWR __dut__._1664_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1595_ __dut__._1767_/A1 __dut__._1593_/X __dut__._1594_/X VGND VGND VPWR
+ VPWR __dut__._1802_/D sky130_fd_sc_hd__a21o_4
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1460__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1094__B1 prod[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1029_ __dut__._1129_/A1 __dut__._1029_/A2 __dut__._1028_/X VGND VGND VPWR
+ VPWR __dut__._1029_/X sky130_fd_sc_hd__a21o_4
XFILLER_9_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1370__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1402_ __dut__.__uuf__._1399_/Y __dut__.__uuf__._1400_/X __dut__.__uuf__._1401_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1402_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1333_ __dut__.__uuf__._1342_/A VGND VGND VPWR VPWR __dut__.__uuf__._1333_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1264_ __dut__.__uuf__._1257_/X __dut__.__uuf__._1254_/X prod[0]
+ prod[1] __dut__.__uuf__._1054_/X VGND VGND VPWR VPWR __dut__._1269_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_100_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1195_ __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR __dut__.__uuf__._1195_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__.__uuf__._1177__A __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1380_ __dut__._1542_/A prod[55] VGND VGND VPWR VPWR __dut__._1380_/X sky130_fd_sc_hd__and2_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__.__uuf__._1091__A3 prod[59] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_190_ _263_/Q _191_/B VGND VGND VPWR VPWR _262_/D sky130_fd_sc_hd__and2_4
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1716_ __dut__._1788_/A __dut__._1833_/Q VGND VGND VPWR VPWR __dut__._1716_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1455__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1087__A __dut__.__uuf__._2008_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1647_ __dut__._1647_/A1 __dut__._1645_/X __dut__._1646_/X VGND VGND VPWR
+ VPWR __dut__._1815_/D sky130_fd_sc_hd__a21o_4
X__dut__._1578_ __dut__._1766_/A __dut__._1797_/Q VGND VGND VPWR VPWR __dut__._1578_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_64_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_13_0___dut__.__uuf__.__clk_source__ clkbuf_3_6_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._2169_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1790__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0___dut__.__uuf__.__clk_source__ __dut__._1411_/X VGND VGND VPWR VPWR clkbuf_0___dut__.__uuf__.__clk_source__/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_174_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1951_ __dut__._1114_/B VGND VGND VPWR VPWR __dut__.__uuf__._1951_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1882_ __dut__.__uuf__._1881_/X __dut__.__uuf__._1880_/B __dut__.__uuf__._1880_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1883_/C sky130_fd_sc_hd__o21ai_4
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._0880_ __dut__._0880_/A __dut__._1856_/Q VGND VGND VPWR VPWR __dut__._0880_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1316_ __dut__.__uuf__._1316_/A VGND VGND VPWR VPWR __dut__.__uuf__._1316_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1501_ rst VGND VGND VPWR VPWR __dut__._1501_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1247_ __dut__.__uuf__._1242_/X __dut__.__uuf__._1239_/X prod[6]
+ prod[7] __dut__.__uuf__._1234_/X VGND VGND VPWR VPWR __dut__._1281_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1178_ __dut__.__uuf__._1236_/A VGND VGND VPWR VPWR __dut__.__uuf__._1189_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1432_ rst VGND VGND VPWR VPWR __dut__._1432_/Y sky130_fd_sc_hd__inv_2
X__dut__._1363_ __dut__._1383_/A1 __dut__._1363_/A2 __dut__._1362_/X VGND VGND VPWR
+ VPWR __dut__._1363_/X sky130_fd_sc_hd__a21o_4
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1294_ __dut__._1324_/A prod[12] VGND VGND VPWR VPWR __dut__._1294_/X sky130_fd_sc_hd__and2_4
XFILLER_42_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_311_ _194_/A _311_/D trst VGND VGND VPWR VPWR _311_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_242_ _242_/A VGND VGND VPWR VPWR _244_/C sky130_fd_sc_hd__inv_2
X_173_ _277_/Q _173_/B VGND VGND VPWR VPWR _276_/D sky130_fd_sc_hd__and2_4
XFILLER_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2074__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__304__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._0903__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2150_ __dut__.__uuf__._2169_/CLK __dut__._1289_/X __dut__.__uuf__._1233_/X
+ VGND VGND VPWR VPWR prod[10] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1101_ __dut__.__uuf__._1093_/X __dut__.__uuf__._1090_/X prod[55]
+ prod[56] __dut__.__uuf__._1100_/X VGND VGND VPWR VPWR __dut__._1379_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_68_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2081_ __dut__.__uuf__._2097_/CLK __dut__._1151_/X __dut__.__uuf__._1546_/X
+ VGND VGND VPWR VPWR __dut__._1152_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1032_ __dut__._1404_/B __dut__.__uuf__._1058_/B VGND VGND VPWR VPWR
+ __dut__.__uuf__._1057_/A sky130_fd_sc_hd__and2_4
XFILLER_68_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1934_ __dut__.__uuf__._1928_/Y __dut__.__uuf__._1929_/Y __dut__.__uuf__._1928_/Y
+ __dut__.__uuf__._1929_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1935_/C sky130_fd_sc_hd__a2bb2o_4
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1865_ __dut__.__uuf__._1862_/Y __dut__.__uuf__._1863_/Y __dut__.__uuf__._1853_/X
+ __dut__.__uuf__._1870_/B VGND VGND VPWR VPWR __dut__.__uuf__._1865_/X sky130_fd_sc_hd__o22a_4
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1796_ __dut__._1058_/B VGND VGND VPWR VPWR __dut__.__uuf__._1796_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._0932_ __dut__._1408_/A __dut__._1882_/Q VGND VGND VPWR VPWR __dut__._0932_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1147__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._0902__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0863_ __dut__._1767_/A1 __dut__._1789_/X __dut__._0862_/X VGND VGND VPWR
+ VPWR __dut__._1851_/D sky130_fd_sc_hd__a21o_4
XFILLER_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1415_ rst VGND VGND VPWR VPWR __dut__._1415_/Y sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_75_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1346_ __dut__._1346_/A prod[38] VGND VGND VPWR VPWR __dut__._1346_/X sky130_fd_sc_hd__and2_4
XFILLER_62_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1277_ __dut__._1277_/A1 __dut__._1277_/A2 __dut__._1276_/X VGND VGND VPWR
+ VPWR __dut__._1277_/X sky130_fd_sc_hd__a21o_4
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_225_ _300_/Q _225_/B VGND VGND VPWR VPWR _299_/D sky130_fd_sc_hd__and2_4
X_156_ _183_/A VGND VGND VPWR VPWR _164_/B sky130_fd_sc_hd__buf_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1689__A2 mp[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_137_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1613__A2 mc[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1650_ __dut__.__uuf__._1654_/A VGND VGND VPWR VPWR __dut__.__uuf__._1650_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1377__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1581_ __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR __dut__.__uuf__._1606_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1129__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2202_ __dut__.__uuf__._2210_/CLK __dut__._1393_/X __dut__.__uuf__._1080_/X
+ VGND VGND VPWR VPWR prod[62] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._2133_ __dut__.__uuf__._2206_/CLK __dut__._1255_/X __dut__.__uuf__._1302_/X
+ VGND VGND VPWR VPWR __dut__._1256_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._2064_ __dut__.__uuf__._2065_/CLK __dut__._1117_/X __dut__.__uuf__._1589_/X
+ VGND VGND VPWR VPWR __dut__._1118_/B sky130_fd_sc_hd__dfrtp_4
X__dut__._1200_ __dut__._1200_/A __dut__._1200_/B VGND VGND VPWR VPWR __dut__._1200_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1272__B prod[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1131_ __dut__._1647_/A1 __dut__._1131_/A2 __dut__._1130_/X VGND VGND VPWR
+ VPWR __dut__._1131_/X sky130_fd_sc_hd__a21o_4
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_108 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1650_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_119 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1140_/A sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1917_ __dut__._1102_/B VGND VGND VPWR VPWR __dut__.__uuf__._1917_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1062_ __dut__._1766_/A __dut__._1062_/B VGND VGND VPWR VPWR __dut__._1062_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA__297__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1848_ __dut__.__uuf__._1859_/A __dut__.__uuf__._1848_/B __dut__.__uuf__._1848_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1850_/B sky130_fd_sc_hd__or3_4
X__dut__.__uuf__._1779_ __dut__.__uuf__._1774_/Y __dut__.__uuf__._1775_/Y __dut__.__uuf__._1776_/X
+ __dut__.__uuf__._1778_/X VGND VGND VPWR VPWR __dut__.__uuf__._1780_/A sky130_fd_sc_hd__a211o_4
XANTENNA___dut__._1851__CLK __dut__._1410_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0915_ __dut__._1383_/A1 prod[54] __dut__._0914_/X VGND VGND VPWR VPWR __dut__._1874_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1728__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1895_ __dut__._1899_/CLK __dut__._1895_/D __dut__._1434_/Y VGND VGND VPWR
+ VPWR __dut__._1895_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1463__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_9_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1258__A3 prod[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1329_ __dut__._1331_/A1 __dut__._1329_/A2 __dut__._1328_/X VGND VGND VPWR
+ VPWR __dut__._1329_/X sky130_fd_sc_hd__a21o_4
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1359__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_208_ _252_/Q _208_/B VGND VGND VPWR VPWR _208_/X sky130_fd_sc_hd__or2_4
X_139_ _238_/B _138_/B _138_/Y _128_/X VGND VGND VPWR VPWR _140_/A sky130_fd_sc_hd__a211o_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2112__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_81_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1733__A __dut__._1609_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1702_ __dut__.__uuf__._1695_/Y __dut__.__uuf__._1696_/Y __dut__.__uuf__._1695_/Y
+ __dut__.__uuf__._1696_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1703_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._1874__CLK __dut__._1917_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1633_ __dut__.__uuf__._1636_/A VGND VGND VPWR VPWR __dut__.__uuf__._1633_/X
+ sky130_fd_sc_hd__buf_2
Xclkbuf_4_0_0_tck clkbuf_4_1_0_tck/A VGND VGND VPWR VPWR _313_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1564_ __dut__.__uuf__._1551_/X __dut__.__uuf__._1547_/X __dut__._1144_/B
+ __dut__.__uuf__._1449_/A __dut__.__uuf__._1563_/X VGND VGND VPWR VPWR __dut__._1143_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1548__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1495_ __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR __dut__.__uuf__._1495_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1680_ __dut__._1788_/A __dut__._1824_/Q VGND VGND VPWR VPWR __dut__._1680_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._2116_ __dut__.__uuf__._2119_/CLK __dut__._1221_/X __dut__.__uuf__._1388_/X
+ VGND VGND VPWR VPWR __dut__._1222_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2047_ __dut__.__uuf__._2049_/CLK __dut__._1083_/X __dut__.__uuf__._1609_/X
+ VGND VGND VPWR VPWR __dut__._1084_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1114_ __dut__._1678_/A __dut__._1114_/B VGND VGND VPWR VPWR __dut__._1114_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1589__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1643__A __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1045_ __dut__._1647_/A1 __dut__._1045_/A2 __dut__._1044_/X VGND VGND VPWR
+ VPWR __dut__._1045_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_38_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1458__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1761__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1878_ __dut__._1919_/CLK __dut__._1878_/D __dut__._1451_/Y VGND VGND VPWR
+ VPWR __dut__._1878_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1897__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1368__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1280_ __dut__._1266_/B VGND VGND VPWR VPWR __dut__.__uuf__._1280_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2158__CLK __dut__.__uuf__._2164_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1616_ __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR __dut__.__uuf__._1616_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1801_ clkbuf_4_6_0_tck/X __dut__._1801_/D __dut__._1528_/Y VGND VGND VPWR
+ VPWR __dut__._1801_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1547_ __dut__.__uuf__._1566_/A VGND VGND VPWR VPWR __dut__.__uuf__._1547_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1732_ __dut__._1788_/A __dut__._1837_/Q VGND VGND VPWR VPWR __dut__._1732_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1478_ __dut__.__uuf__._1466_/X __dut__.__uuf__._1462_/X __dut__._1186_/B
+ __dut__.__uuf__._1471_/X __dut__.__uuf__._1477_/X VGND VGND VPWR VPWR __dut__._1185_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._0910__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1663_ __dut__._1767_/A1 __dut__._1661_/X __dut__._1662_/X VGND VGND VPWR
+ VPWR __dut__._1819_/D sky130_fd_sc_hd__a21o_4
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1594_ __dut__._1766_/A __dut__._1800_/Q VGND VGND VPWR VPWR __dut__._1594_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_17_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_7_0_tck clkbuf_3_7_0_tck/A VGND VGND VPWR VPWR clkbuf_3_7_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1028_ __dut__._1078_/A __dut__._1028_/B VGND VGND VPWR VPWR __dut__._1028_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1725__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1401_ __dut__.__uuf__._1401_/A VGND VGND VPWR VPWR __dut__.__uuf__._1401_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1912__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1332_ __dut__.__uuf__._1329_/X __dut__.__uuf__._1331_/X __dut__._1246_/B
+ __dut__.__uuf__._1329_/X VGND VGND VPWR VPWR __dut__._1245_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1263_ __dut__.__uuf__._1263_/A VGND VGND VPWR VPWR __dut__.__uuf__._1263_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_98_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1194_ __dut__.__uuf__._1204_/A VGND VGND VPWR VPWR __dut__.__uuf__._1194_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_27_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1715_ __dut__._1719_/A1 __dut__._1713_/X __dut__._1714_/X VGND VGND VPWR
+ VPWR __dut__._1832_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1736__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1646_ __dut__._1646_/A __dut__._1814_/Q VGND VGND VPWR VPWR __dut__._1646_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_77_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1577_ __dut__._1543_/Y mc[17] __dut__._1576_/X VGND VGND VPWR VPWR __dut__._1577_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1471__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0___dut__.__uuf__.__clk_source__ clkbuf_3_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_5_0___dut__.__uuf__.__clk_source__/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_167_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1950_ __dut__.__uuf__._1990_/A __dut__.__uuf__._1950_/B __dut__.__uuf__._1950_/C
+ VGND VGND VPWR VPWR __dut__._1107_/A2 sky130_fd_sc_hd__and3_4
X__dut__.__uuf__._1881_ __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR __dut__.__uuf__._1881_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__284__CLK _290_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1315_ __dut__.__uuf__._1303_/X __dut__.__uuf__._1313_/X __dut__._1252_/B
+ __dut__.__uuf__._1314_/X VGND VGND VPWR VPWR __dut__._1251_/A2 sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._1556__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1500_ rst VGND VGND VPWR VPWR __dut__._1500_/Y sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1246_ __dut__.__uuf__._1248_/A VGND VGND VPWR VPWR __dut__.__uuf__._1246_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1177_ __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR __dut__.__uuf__._1236_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1431_ rst VGND VGND VPWR VPWR __dut__._1431_/Y sky130_fd_sc_hd__inv_2
X__dut__._1362_ __dut__._1378_/A prod[46] VGND VGND VPWR VPWR __dut__._1362_/X sky130_fd_sc_hd__and2_4
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1808__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1293_ __dut__._1293_/A1 __dut__._1293_/A2 __dut__._1292_/X VGND VGND VPWR
+ VPWR __dut__._1293_/X sky130_fd_sc_hd__a21o_4
X_310_ _314_/CLK _310_/D trst VGND VGND VPWR VPWR _310_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_241_ tms _240_/X _128_/X VGND VGND VPWR VPWR _306_/D sky130_fd_sc_hd__a21o_4
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_20_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_172_ _278_/Q _172_/B VGND VGND VPWR VPWR _277_/D sky130_fd_sc_hd__or2_4
XFILLER_6_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1466__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1629_ __dut__._1543_/Y mc[29] __dut__._1628_/X VGND VGND VPWR VPWR __dut__._1629_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_92_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1376__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1100_ __dut__.__uuf__._1100_/A VGND VGND VPWR VPWR __dut__.__uuf__._1100_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2080_ __dut__.__uuf__._2097_/CLK __dut__._1149_/X __dut__.__uuf__._1550_/X
+ VGND VGND VPWR VPWR __dut__._1150_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1031_ __dut__.__uuf__._1031_/A VGND VGND VPWR VPWR __dut__.__uuf__._1058_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1933_ __dut__.__uuf__._1933_/A VGND VGND VPWR VPWR __dut__._1105_/A2
+ sky130_fd_sc_hd__inv_2
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1864_ __dut__._1557_/X VGND VGND VPWR VPWR __dut__.__uuf__._1870_/B
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1795_ __dut__.__uuf__._1828_/A __dut__.__uuf__._1795_/B __dut__.__uuf__._1795_/C
+ VGND VGND VPWR VPWR __dut__._1051_/A2 sky130_fd_sc_hd__and3_4
X__dut__._0931_ __dut__._1395_/A1 prod[62] __dut__._0930_/X VGND VGND VPWR VPWR __dut__._1882_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._0862_ __dut__._1766_/A __dut__._1845_/Q VGND VGND VPWR VPWR __dut__._0862_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1286__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1229_ __dut__.__uuf__._1233_/A VGND VGND VPWR VPWR __dut__.__uuf__._1229_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_74_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1414_ rst VGND VGND VPWR VPWR __dut__._1414_/Y sky130_fd_sc_hd__inv_2
X__dut__._1345_ __dut__._1349_/A1 __dut__._1345_/A2 __dut__._1344_/X VGND VGND VPWR
+ VPWR __dut__._1345_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_68_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1083__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1276_ __dut__._1276_/A prod[3] VGND VGND VPWR VPWR __dut__._1276_/X sky130_fd_sc_hd__and2_4
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_224_ _301_/Q _299_/Q _232_/A VGND VGND VPWR VPWR _298_/D sky130_fd_sc_hd__o21a_4
X_155_ _193_/B VGND VGND VPWR VPWR _183_/A sky130_fd_sc_hd__inv_2
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0897__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1556__A __dut__.__uuf__._1720_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1580_ __dut__.__uuf__._1580_/A VGND VGND VPWR VPWR __dut__.__uuf__._1580_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2201_ __dut__.__uuf__._2210_/CLK __dut__._1391_/X __dut__.__uuf__._1082_/X
+ VGND VGND VPWR VPWR prod[61] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2132_ __dut__.__uuf__._2206_/CLK __dut__._1253_/X __dut__.__uuf__._1307_/X
+ VGND VGND VPWR VPWR __dut__._1254_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2063_ __dut__.__uuf__._2065_/CLK __dut__._1115_/X __dut__.__uuf__._1590_/X
+ VGND VGND VPWR VPWR __dut__._1116_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1130_ __dut__._1130_/A __dut__._1130_/B VGND VGND VPWR VPWR __dut__._1130_/X
+ sky130_fd_sc_hd__and2_4
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpsn_inst_psn_buff_109 __dut__._1678_/A VGND VGND VPWR VPWR __dut__._1646_/A sky130_fd_sc_hd__buf_2
XFILLER_12_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1916_ __dut__.__uuf__._1938_/A __dut__.__uuf__._1916_/B __dut__.__uuf__._1916_/C
+ VGND VGND VPWR VPWR __dut__._1095_/A2 sky130_fd_sc_hd__and3_4
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1061_ __dut__._1071_/A1 __dut__._1061_/A2 __dut__._1060_/X VGND VGND VPWR
+ VPWR __dut__._1061_/X sky130_fd_sc_hd__a21o_4
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1847_ __dut__.__uuf__._1841_/Y __dut__.__uuf__._1842_/Y __dut__.__uuf__._1841_/Y
+ __dut__.__uuf__._1842_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1848_/C sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1778_ __dut__.__uuf__._1774_/Y __dut__.__uuf__._1775_/Y __dut__.__uuf__._1743_/X
+ __dut__.__uuf__._1783_/B VGND VGND VPWR VPWR __dut__.__uuf__._1778_/X sky130_fd_sc_hd__o22a_4
X__dut__._0914_ __dut__._1378_/A __dut__._1873_/Q VGND VGND VPWR VPWR __dut__._0914_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1894_ __dut__._1899_/CLK __dut__._1894_/D __dut__._1435_/Y VGND VGND VPWR
+ VPWR __dut__._1894_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1744__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1328_ __dut__._1378_/A prod[29] VGND VGND VPWR VPWR __dut__._1328_/X sky130_fd_sc_hd__and2_4
XFILLER_15_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1259_ __dut__._1787_/A1 __dut__._1259_/A2 __dut__._1258_/X VGND VGND VPWR
+ VPWR __dut__._1259_/X sky130_fd_sc_hd__a21o_4
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_207_ _211_/A VGND VGND VPWR VPWR _208_/B sky130_fd_sc_hd__inv_2
X_138_ _307_/Q _138_/B VGND VGND VPWR VPWR _138_/Y sky130_fd_sc_hd__nor2_4
XFILLER_97_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1654__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1701_ __dut__.__uuf__._1868_/A VGND VGND VPWR VPWR __dut__.__uuf__._1749_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1632_ __dut__.__uuf__._1636_/A VGND VGND VPWR VPWR __dut__.__uuf__._1632_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1563_ __dut__._1649_/X __dut__.__uuf__._1078_/A __dut__._1146_/B
+ __dut__.__uuf__._1660_/A VGND VGND VPWR VPWR __dut__.__uuf__._1563_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1494_ __dut__.__uuf__._1536_/A VGND VGND VPWR VPWR __dut__.__uuf__._1494_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_88_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1564__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2115_ __dut__.__uuf__._2138_/CLK __dut__._1219_/X __dut__.__uuf__._1393_/X
+ VGND VGND VPWR VPWR __dut__._1220_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2046_ __dut__.__uuf__._2049_/CLK __dut__._1081_/X __dut__.__uuf__._1610_/X
+ VGND VGND VPWR VPWR __dut__._1082_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0908__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1113_ __dut__._1129_/A1 __dut__._1113_/A2 __dut__._1112_/X VGND VGND VPWR
+ VPWR __dut__._1113_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1589__A2 mc[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1044_ __dut__._1044_/A __dut__._1044_/B VGND VGND VPWR VPWR __dut__._1044_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1761__A2 mp[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1877_ __dut__._1919_/CLK __dut__._1877_/D __dut__._1452_/Y VGND VGND VPWR
+ VPWR __dut__._1877_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1474__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1029__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1384__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1841__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1615_ __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR __dut__.__uuf__._1615_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1800_ __dut__._1410_/B __dut__._1800_/D __dut__._1529_/Y VGND VGND VPWR
+ VPWR __dut__._1800_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1546_ __dut__.__uuf__._1550_/A VGND VGND VPWR VPWR __dut__.__uuf__._1546_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_1_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1731_ __dut__._1731_/A1 __dut__._1729_/X __dut__._1730_/X VGND VGND VPWR
+ VPWR __dut__._1836_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1477_ __dut__._1741_/X __dut__.__uuf__._1472_/X __dut__._1188_/B
+ __dut__.__uuf__._1473_/X VGND VGND VPWR VPWR __dut__.__uuf__._1477_/X sky130_fd_sc_hd__o22a_4
XANTENNA___dut__.__uuf__._1919__A __dut__._0865_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1662_ __dut__._1766_/A __dut__._1818_/Q VGND VGND VPWR VPWR __dut__._1662_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1593_ __dut__._1543_/Y mc[20] __dut__._1592_/X VGND VGND VPWR VPWR __dut__._1593_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1259__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2029_ __dut__.__uuf__._2083_/CLK __dut__._1047_/X __dut__.__uuf__._1632_/X
+ VGND VGND VPWR VPWR __dut__._1048_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_50_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2102__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_71_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1027_ __dut__._1129_/A1 __dut__._1027_/A2 __dut__._1026_/X VGND VGND VPWR
+ VPWR __dut__._1027_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1469__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1864__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_112_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1725__A2 mp[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1400_ __dut__.__uuf__._1400_/A VGND VGND VPWR VPWR __dut__.__uuf__._1400_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1331_ __dut__.__uuf__._1330_/Y __dut__.__uuf__._1323_/X __dut__.__uuf__._1324_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1331_/X sky130_fd_sc_hd__o21a_4
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1262_ __dut__.__uuf__._1257_/X __dut__.__uuf__._1254_/X prod[1]
+ prod[2] __dut__.__uuf__._1249_/X VGND VGND VPWR VPWR __dut__._1271_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1193_ __dut__.__uuf__._1236_/A VGND VGND VPWR VPWR __dut__.__uuf__._1204_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_100_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1661__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1529_ __dut__.__uuf__._1529_/A VGND VGND VPWR VPWR __dut__.__uuf__._1529_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_89_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1649__A __dut__.__uuf__._1649_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1714_ __dut__._1766_/A __dut__._1831_/Q VGND VGND VPWR VPWR __dut__._1714_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_98_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1645_ __dut__._1543_/Y mp[0] __dut__._1644_/X VGND VGND VPWR VPWR __dut__._1645_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1576_ __dut__._1788_/A __dut__._1798_/Q VGND VGND VPWR VPWR __dut__._1576_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1752__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1662__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1643__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1880_ __dut__.__uuf__._1914_/A __dut__.__uuf__._1880_/B __dut__.__uuf__._1880_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1883_/B sky130_fd_sc_hd__or3_4
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2007__A1 done VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1314_ __dut__.__uuf__._1314_/A VGND VGND VPWR VPWR __dut__.__uuf__._1314_/X
+ sky130_fd_sc_hd__buf_2
Xclkbuf_3_6_0_tck clkbuf_3_7_0_tck/A VGND VGND VPWR VPWR clkbuf_3_6_0_tck/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1245_ __dut__.__uuf__._1242_/X __dut__.__uuf__._1239_/X prod[7]
+ prod[8] __dut__.__uuf__._1234_/X VGND VGND VPWR VPWR __dut__._1283_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1176_ __dut__.__uuf__._1168_/X __dut__.__uuf__._1165_/X prod[30]
+ prod[31] __dut__.__uuf__._1175_/X VGND VGND VPWR VPWR __dut__._1329_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1430_ rst VGND VGND VPWR VPWR __dut__._1430_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1361_ __dut__._1383_/A1 __dut__._1361_/A2 __dut__._1360_/X VGND VGND VPWR
+ VPWR __dut__._1361_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1572__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1292_ __dut__._1324_/A prod[11] VGND VGND VPWR VPWR __dut__._1292_/X sky130_fd_sc_hd__and2_4
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0916__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_240_ _297_/Q _306_/Q VGND VGND VPWR VPWR _240_/X sky130_fd_sc_hd__or2_4
XFILLER_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_171_ _279_/Q _173_/B VGND VGND VPWR VPWR _278_/D sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_13_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1628_ __dut__._1788_/A __dut__._1811_/Q VGND VGND VPWR VPWR __dut__._1628_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1482__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1559_ __dut__._1767_/A1 __dut__._1557_/X __dut__._1558_/X VGND VGND VPWR
+ VPWR __dut__._1793_/D sky130_fd_sc_hd__a21o_4
XFILLER_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1625__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2003__A __dut__.__uuf__._2003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1902__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1030_ __dut__.__uuf__._1061_/A __dut__.__uuf__._1061_/B VGND VGND
+ VPWR VPWR __dut__.__uuf__._1031_/A sky130_fd_sc_hd__or2_4
XANTENNA___dut__._1392__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__313__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1932_ __dut__.__uuf__._1928_/Y __dut__.__uuf__._1929_/Y __dut__.__uuf__._1886_/X
+ __dut__.__uuf__._1931_/X VGND VGND VPWR VPWR __dut__.__uuf__._1933_/A sky130_fd_sc_hd__a211o_4
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1863_ __dut__._1076_/B VGND VGND VPWR VPWR __dut__.__uuf__._1863_/Y
+ sky130_fd_sc_hd__inv_2
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1794_ __dut__.__uuf__._1771_/X __dut__.__uuf__._1793_/B __dut__.__uuf__._1793_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1795_/C sky130_fd_sc_hd__o21ai_4
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0930_ __dut__._1542_/A __dut__._1881_/Q VGND VGND VPWR VPWR __dut__._0930_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1228_ __dut__.__uuf__._1227_/X __dut__.__uuf__._1223_/X prod[13]
+ prod[14] __dut__.__uuf__._1219_/X VGND VGND VPWR VPWR __dut__._1295_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1413_ rst VGND VGND VPWR VPWR __dut__._1413_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1159_ __dut__.__uuf__._1159_/A VGND VGND VPWR VPWR __dut__.__uuf__._1159_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1344_ __dut__._1344_/A prod[37] VGND VGND VPWR VPWR __dut__._1344_/X sky130_fd_sc_hd__and2_4
XFILLER_74_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1607__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1275_ __dut__._1275_/A1 __dut__._1275_/A2 __dut__._1274_/X VGND VGND VPWR
+ VPWR __dut__._1275_/X sky130_fd_sc_hd__a21o_4
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_223_ _304_/Q _225_/B VGND VGND VPWR VPWR _297_/D sky130_fd_sc_hd__and2_4
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_154_ _238_/A _311_/Q _154_/C _242_/A VGND VGND VPWR VPWR _193_/B sky130_fd_sc_hd__or4_4
XANTENNA___dut__._1477__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__274__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._2200_ __dut__.__uuf__._2200_/CLK __dut__._1389_/X __dut__.__uuf__._1084_/X
+ VGND VGND VPWR VPWR prod[60] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2131_ __dut__.__uuf__._2206_/CLK __dut__._1251_/X __dut__.__uuf__._1311_/X
+ VGND VGND VPWR VPWR __dut__._1252_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2062_ __dut__.__uuf__._2065_/CLK __dut__._1113_/X __dut__.__uuf__._1591_/X
+ VGND VGND VPWR VPWR __dut__._1114_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1915_ __dut__.__uuf__._1881_/X __dut__.__uuf__._1914_/B __dut__.__uuf__._1914_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1916_/C sky130_fd_sc_hd__o21ai_4
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1060_ __dut__._1074_/A __dut__._1060_/B VGND VGND VPWR VPWR __dut__._1060_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1846_ __dut__.__uuf__._1846_/A VGND VGND VPWR VPWR __dut__._1073_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1777_ __dut__._1593_/X VGND VGND VPWR VPWR __dut__.__uuf__._1783_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_20_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._0913_ __dut__._1383_/A1 prod[53] __dut__._0912_/X VGND VGND VPWR VPWR __dut__._1873_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1893_ __dut__._1899_/CLK __dut__._1893_/D __dut__._1436_/Y VGND VGND VPWR
+ VPWR __dut__._1893_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_80_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2209__CLK __dut__.__uuf__._2210_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_74_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1327_ __dut__._1327_/A1 __dut__._1327_/A2 __dut__._1326_/X VGND VGND VPWR
+ VPWR __dut__._1327_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1760__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1258_ __dut__._1786_/A __dut__._1258_/B VGND VGND VPWR VPWR __dut__._1258_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1189_ __dut__._1193_/A1 __dut__._1189_/A2 __dut__._1188_/X VGND VGND VPWR
+ VPWR __dut__._1189_/X sky130_fd_sc_hd__a21o_4
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_206_ _206_/A _250_/Q _249_/Q VGND VGND VPWR VPWR _211_/A sky130_fd_sc_hd__or3_4
X_137_ _311_/Q VGND VGND VPWR VPWR _238_/B sky130_fd_sc_hd__inv_2
XFILLER_99_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__._1000__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_142_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1670__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1700_ __dut__.__uuf__._1700_/A VGND VGND VPWR VPWR __dut__._1021_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1631_ __dut__.__uuf__._1637_/A VGND VGND VPWR VPWR __dut__.__uuf__._1636_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1562_ __dut__.__uuf__._1569_/A VGND VGND VPWR VPWR __dut__.__uuf__._1562_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1493_ __dut__.__uuf__._1535_/A VGND VGND VPWR VPWR __dut__.__uuf__._1493_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._2114_ __dut__.__uuf__._2114_/CLK __dut__._1217_/X __dut__.__uuf__._1398_/X
+ VGND VGND VPWR VPWR __dut__._1218_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2045_ __dut__.__uuf__._2049_/CLK __dut__._1079_/X __dut__.__uuf__._1611_/X
+ VGND VGND VPWR VPWR __dut__._1080_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_29_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1580__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1112_ __dut__._1112_/A __dut__._1112_/B VGND VGND VPWR VPWR __dut__._1112_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1043_ __dut__._1647_/A1 __dut__._1043_/A2 __dut__._1042_/X VGND VGND VPWR
+ VPWR __dut__._1043_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1829_ __dut__._1070_/B VGND VGND VPWR VPWR __dut__.__uuf__._1829_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._0924__A __dut__._1542_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1876_ __dut__._1919_/CLK __dut__._1876_/D __dut__._1453_/Y VGND VGND VPWR
+ VPWR __dut__._1876_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__312__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1490__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1793__CLK __dut__._1410_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1614_ __dut__.__uuf__._1618_/A VGND VGND VPWR VPWR __dut__.__uuf__._1614_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1545_ __dut__.__uuf__._1530_/X __dut__.__uuf__._1526_/X __dut__._1154_/B
+ __dut__.__uuf__._1535_/X __dut__.__uuf__._1544_/X VGND VGND VPWR VPWR __dut__._1153_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1260__B1 prod[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1730_ __dut__._1766_/A __dut__._1835_/Q VGND VGND VPWR VPWR __dut__._1730_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1476_ __dut__.__uuf__._1486_/A VGND VGND VPWR VPWR __dut__.__uuf__._1476_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1661_ __dut__._1543_/Y mp[4] __dut__._1660_/X VGND VGND VPWR VPWR __dut__._1661_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__._1592_ __dut__._1788_/A __dut__._1802_/Q VGND VGND VPWR VPWR __dut__._1592_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2028_ __dut__.__uuf__._2083_/CLK __dut__._1045_/X __dut__.__uuf__._1633_/X
+ VGND VGND VPWR VPWR __dut__._1046_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._1079__B1 __dut__._1132_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_psn_inst_psn_buff_43_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1026_ __dut__._1128_/A __dut__._1026_/B VGND VGND VPWR VPWR __dut__._1026_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_40_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1485__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1859_ __dut__._1883_/CLK __dut__._1859_/D __dut__._1470_/Y VGND VGND VPWR
+ VPWR __dut__._1859_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_105_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2077__CLK __dut__.__uuf__._2107_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1330_ __dut__._1248_/B VGND VGND VPWR VPWR __dut__.__uuf__._1330_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1261_ __dut__.__uuf__._1263_/A VGND VGND VPWR VPWR __dut__.__uuf__._1261_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1192_ __dut__.__uuf__._1183_/X __dut__.__uuf__._1180_/X prod[25]
+ prod[26] __dut__.__uuf__._1191_/X VGND VGND VPWR VPWR __dut__._1319_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1661__A2 mp[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__.__uuf__._1490__A __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1177__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1528_ __dut__.__uuf__._1509_/X __dut__.__uuf__._1526_/X __dut__._1162_/B
+ __dut__.__uuf__._1514_/X __dut__.__uuf__._1527_/X VGND VGND VPWR VPWR __dut__._1161_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1713_ __dut__._1543_/Y mp[16] __dut__._1712_/X VGND VGND VPWR VPWR __dut__._1713_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1459_ __dut__._1757_/X __dut__.__uuf__._1451_/X __dut__._1196_/B
+ __dut__.__uuf__._1452_/X VGND VGND VPWR VPWR __dut__.__uuf__._1459_/X sky130_fd_sc_hd__o22a_4
XFILLER_89_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1644_ __dut__._1788_/A __dut__._1815_/Q VGND VGND VPWR VPWR __dut__._1644_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_49_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1575_ __dut__._1767_/A1 __dut__._1573_/X __dut__._1574_/X VGND VGND VPWR
+ VPWR __dut__._1797_/D sky130_fd_sc_hd__a21o_4
XFILLER_66_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1101__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1009_ __dut__._1129_/A1 __dut__._1009_/A2 __dut__._1008_/X VGND VGND VPWR
+ VPWR __dut__._1009_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._0915__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1831__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__194__A _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1313_ __dut__.__uuf__._1312_/Y __dut__.__uuf__._1297_/X __dut__.__uuf__._1299_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1313_/X sky130_fd_sc_hd__o21a_4
X__dut__.__uuf__._1244_ __dut__.__uuf__._1248_/A VGND VGND VPWR VPWR __dut__.__uuf__._1244_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1175_ __dut__.__uuf__._1175_/A VGND VGND VPWR VPWR __dut__.__uuf__._1175_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_59_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1360_ __dut__._1378_/A prod[45] VGND VGND VPWR VPWR __dut__._1360_/X sky130_fd_sc_hd__and2_4
XFILLER_74_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1291_ __dut__._1291_/A1 __dut__._1291_/A2 __dut__._1290_/X VGND VGND VPWR
+ VPWR __dut__._1291_/X sky130_fd_sc_hd__a21o_4
XFILLER_82_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_tck_A tck VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_170_ _280_/Q _172_/B VGND VGND VPWR VPWR _279_/D sky130_fd_sc_hd__or2_4
XFILLER_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1854__CLK clkbuf_4_5_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1627_ __dut__._1647_/A1 __dut__._1625_/X __dut__._1626_/X VGND VGND VPWR
+ VPWR __dut__._1810_/D sky130_fd_sc_hd__a21o_4
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1558_ __dut__._1766_/A __dut__._1792_/Q VGND VGND VPWR VPWR __dut__._1558_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1625__A2 mc[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1489_ rst VGND VGND VPWR VPWR __dut__._1489_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_299_ _194_/A _299_/D trst VGND VGND VPWR VPWR _299_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1561__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_psn_inst_psn_buff_172_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1392__B prod[61] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1931_ __dut__.__uuf__._1928_/Y __dut__.__uuf__._1929_/Y __dut__.__uuf__._1908_/X
+ __dut__.__uuf__._1935_/B VGND VGND VPWR VPWR __dut__.__uuf__._1931_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1862_ __dut__._1082_/B VGND VGND VPWR VPWR __dut__.__uuf__._1862_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1877__CLK __dut__._1919_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1793_ __dut__.__uuf__._1804_/A __dut__.__uuf__._1793_/B __dut__.__uuf__._1793_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1795_/B sky130_fd_sc_hd__or3_4
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1227_ __dut__.__uuf__._1466_/A VGND VGND VPWR VPWR __dut__.__uuf__._1227_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1158_ __dut__.__uuf__._1153_/X __dut__.__uuf__._1149_/X prod[36]
+ prod[37] __dut__.__uuf__._1145_/X VGND VGND VPWR VPWR __dut__._1341_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1412_ rst VGND VGND VPWR VPWR __dut__._1412_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1343_ __dut__._1343_/A1 __dut__._1343_/A2 __dut__._1342_/X VGND VGND VPWR
+ VPWR __dut__._1343_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1089_ __dut__.__uuf__._1450_/A VGND VGND VPWR VPWR __dut__.__uuf__._1149_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1274_ __dut__._1274_/A prod[2] VGND VGND VPWR VPWR __dut__._1274_/X sky130_fd_sc_hd__and2_4
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_222_ _222_/A _297_/Q VGND VGND VPWR VPWR _296_/D sky130_fd_sc_hd__and2_4
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_153_ _314_/Q _313_/Q VGND VGND VPWR VPWR _242_/A sky130_fd_sc_hd__or2_4
XANTENNA___dut__._1758__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0989_ __dut__._0989_/A1 prod[26] __dut__._0988_/X VGND VGND VPWR VPWR __dut__._1911_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_78_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1493__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_tck clkbuf_3_5_0_tck/A VGND VGND VPWR VPWR clkbuf_3_5_0_tck/X sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1668__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2130_ __dut__.__uuf__._2206_/CLK __dut__._1249_/X __dut__.__uuf__._1316_/X
+ VGND VGND VPWR VPWR __dut__._1250_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2061_ __dut__.__uuf__._2065_/CLK __dut__._1111_/X __dut__.__uuf__._1592_/X
+ VGND VGND VPWR VPWR __dut__._1112_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_96_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1914_ __dut__.__uuf__._1914_/A __dut__.__uuf__._1914_/B __dut__.__uuf__._1914_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1916_/B sky130_fd_sc_hd__or3_4
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1845_ __dut__.__uuf__._1841_/Y __dut__.__uuf__._1842_/Y __dut__.__uuf__._1831_/X
+ __dut__.__uuf__._1844_/X VGND VGND VPWR VPWR __dut__.__uuf__._1846_/A sky130_fd_sc_hd__a211o_4
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1776_ __dut__.__uuf__._1941_/A VGND VGND VPWR VPWR __dut__.__uuf__._1776_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1578__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1773__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0912_ __dut__._1378_/A __dut__._1872_/Q VGND VGND VPWR VPWR __dut__._0912_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1892_ __dut__._1902_/CLK __dut__._1892_/D __dut__._1437_/Y VGND VGND VPWR
+ VPWR __dut__._1892_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_73_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1326_ __dut__._1378_/A prod[28] VGND VGND VPWR VPWR __dut__._1326_/X sky130_fd_sc_hd__and2_4
XFILLER_43_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1257_ __dut__._1787_/A1 __dut__._1257_/A2 __dut__._1256_/X VGND VGND VPWR
+ VPWR __dut__._1257_/X sky130_fd_sc_hd__a21o_4
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1188_ __dut__._1188_/A __dut__._1188_/B VGND VGND VPWR VPWR __dut__._1188_/X
+ sky130_fd_sc_hd__and2_4
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_205_ _248_/Q VGND VGND VPWR VPWR _206_/A sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1488__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_136_ _312_/Q _138_/B _135_/X _128_/X VGND VGND VPWR VPWR _312_/D sky130_fd_sc_hd__a211o_4
XFILLER_99_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_135_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1630_ __dut__.__uuf__._1630_/A VGND VGND VPWR VPWR __dut__.__uuf__._1630_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1561_ __dut__.__uuf__._1551_/X __dut__.__uuf__._1547_/X __dut__._1146_/B
+ __dut__.__uuf__._1449_/A __dut__.__uuf__._1560_/X VGND VGND VPWR VPWR __dut__._1145_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1915__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1492_ __dut__.__uuf__._1508_/A VGND VGND VPWR VPWR __dut__.__uuf__._1492_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2113_ __dut__.__uuf__._2114_/CLK __dut__._1215_/X __dut__.__uuf__._1404_/X
+ VGND VGND VPWR VPWR __dut__._1216_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2044_ __dut__.__uuf__._2049_/CLK __dut__._1077_/X __dut__.__uuf__._1614_/X
+ VGND VGND VPWR VPWR __dut__._1078_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__241__A1 tms VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1111_ __dut__._1129_/A1 __dut__._1111_/A2 __dut__._1110_/X VGND VGND VPWR
+ VPWR __dut__._1111_/X sky130_fd_sc_hd__a21o_4
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1042_ __dut__._1042_/A __dut__._1042_/B VGND VGND VPWR VPWR __dut__._1042_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1828_ __dut__.__uuf__._1828_/A __dut__.__uuf__._1828_/B __dut__.__uuf__._1828_/C
+ VGND VGND VPWR VPWR __dut__._1063_/A2 sky130_fd_sc_hd__and3_4
X__dut__.__uuf__._1759_ __dut__.__uuf__._1752_/Y __dut__.__uuf__._1753_/Y __dut__.__uuf__._1752_/Y
+ __dut__.__uuf__._1753_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1760_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1875_ __dut__._1883_/CLK __dut__._1875_/D __dut__._1454_/Y VGND VGND VPWR
+ VPWR __dut__._1875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_7_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1309_ __dut__._1319_/A1 __dut__._1309_/A2 __dut__._1308_/X VGND VGND VPWR
+ VPWR __dut__._1309_/X sky130_fd_sc_hd__a21o_4
XFILLER_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1737__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0___dut__.__uuf__.__clk_source__ clkbuf_4_9_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2138_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_100_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0___dut__.__uuf__.__clk_source__ clkbuf_0___dut__.__uuf__.__clk_source__/X
+ VGND VGND VPWR VPWR clkbuf_2_1_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__287__CLK _314_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1613_ __dut__.__uuf__._1637_/A VGND VGND VPWR VPWR __dut__.__uuf__._1618_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1544_ __dut__._1669_/X __dut__.__uuf__._1536_/X __dut__._1156_/B
+ __dut__.__uuf__._1537_/X VGND VGND VPWR VPWR __dut__.__uuf__._1544_/X sky130_fd_sc_hd__o22a_4
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1475_ __dut__.__uuf__._1466_/X __dut__.__uuf__._1462_/X __dut__._1188_/B
+ __dut__.__uuf__._1471_/X __dut__.__uuf__._1474_/X VGND VGND VPWR VPWR __dut__._1187_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1660_ __dut__._1788_/A __dut__._1819_/Q VGND VGND VPWR VPWR __dut__._1660_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1591_ __dut__._1647_/A1 __dut__._1589_/X __dut__._1590_/X VGND VGND VPWR
+ VPWR __dut__._1801_/D sky130_fd_sc_hd__a21o_4
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2027_ __dut__.__uuf__._2043_/CLK __dut__._1043_/X __dut__.__uuf__._1634_/X
+ VGND VGND VPWR VPWR __dut__._1044_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._1079__B2 __dut__.__uuf__._1069_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_36_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1025_ __dut__._1129_/A1 __dut__._1025_/A2 __dut__._1024_/X VGND VGND VPWR
+ VPWR __dut__._1025_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1766__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1858_ __dut__._1883_/CLK __dut__._1858_/D __dut__._1471_/Y VGND VGND VPWR
+ VPWR __dut__._1858_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1789_ __dut__._1543_/Y mc[6] __dut__._1788_/X VGND VGND VPWR VPWR __dut__._1789_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_0_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1006__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._0933__A2 prod[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1676__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__307__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1260_ __dut__.__uuf__._1257_/X __dut__.__uuf__._1254_/X prod[2]
+ prod[3] __dut__.__uuf__._1249_/X VGND VGND VPWR VPWR __dut__._1273_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1191_ __dut__.__uuf__._1249_/A VGND VGND VPWR VPWR __dut__.__uuf__._1191_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_3_0_tck_A clkbuf_2_3_0_tck/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__.__uuf__._2021__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1586__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1527_ __dut__._1689_/X __dut__.__uuf__._1515_/X __dut__._1164_/B
+ __dut__.__uuf__._1516_/X VGND VGND VPWR VPWR __dut__.__uuf__._1527_/X sky130_fd_sc_hd__o22a_4
XANTENNA__302__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1712_ __dut__._1788_/A __dut__._1832_/Q VGND VGND VPWR VPWR __dut__._1712_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1458_ __dut__.__uuf__._1465_/A VGND VGND VPWR VPWR __dut__.__uuf__._1458_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_89_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1643_ __dut__._1647_/A1 __dut__._1641_/X __dut__._1642_/X VGND VGND VPWR
+ VPWR __dut__._1814_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1389_ __dut__._1224_/B VGND VGND VPWR VPWR __dut__.__uuf__._1389_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA___dut__.__uuf__._1946__A __dut__.__uuf__._1946_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1574_ __dut__._1766_/A __dut__._1796_/Q VGND VGND VPWR VPWR __dut__._1574_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1008_ __dut__._1008_/A __dut__._1008_/B VGND VGND VPWR VPWR __dut__._1008_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1496__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2044__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1312_ __dut__._1254_/B VGND VGND VPWR VPWR __dut__.__uuf__._1312_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1243_ __dut__.__uuf__._1242_/X __dut__.__uuf__._1239_/X prod[8]
+ prod[9] __dut__.__uuf__._1234_/X VGND VGND VPWR VPWR __dut__._1285_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_86_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1174_ __dut__.__uuf__._1174_/A VGND VGND VPWR VPWR __dut__.__uuf__._1174_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1095__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1290_ __dut__._1770_/A prod[10] VGND VGND VPWR VPWR __dut__._1290_/X sky130_fd_sc_hd__and2_4
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1626_ __dut__._1626_/A __dut__._1809_/Q VGND VGND VPWR VPWR __dut__._1626_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1557_ __dut__._1543_/Y mc[12] __dut__._1556_/X VGND VGND VPWR VPWR __dut__._1557_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_65_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2067__CLK __dut__.__uuf__._2119_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1488_ rst VGND VGND VPWR VPWR __dut__._1488_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_298_ _306_/CLK _298_/D trst VGND VGND VPWR VPWR _298_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1561__A2 mc[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_165_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1077__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1930_ __dut__._1789_/X VGND VGND VPWR VPWR __dut__.__uuf__._1935_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_64_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1861_ __dut__.__uuf__._1883_/A __dut__.__uuf__._1861_/B __dut__.__uuf__._1861_/C
+ VGND VGND VPWR VPWR __dut__._1075_/A2 sky130_fd_sc_hd__and3_4
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1792_ __dut__.__uuf__._1786_/Y __dut__.__uuf__._1787_/Y __dut__.__uuf__._1786_/Y
+ __dut__.__uuf__._1787_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1793_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1226_ __dut__.__uuf__._1226_/A VGND VGND VPWR VPWR __dut__.__uuf__._1466_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_59_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1157_ __dut__.__uuf__._1159_/A VGND VGND VPWR VPWR __dut__.__uuf__._1157_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1411_ __dut__._1543_/Y clk __dut__._1410_/X VGND VGND VPWR VPWR __dut__._1411_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA_clkbuf_1_0_0_tck_A clkbuf_0_tck/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1088_ __dut__.__uuf__._1099_/A VGND VGND VPWR VPWR __dut__.__uuf__._1088_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1342_ __dut__._1342_/A prod[36] VGND VGND VPWR VPWR __dut__._1342_/X sky130_fd_sc_hd__and2_4
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1273_ __dut__._1273_/A1 __dut__._1273_/A2 __dut__._1272_/X VGND VGND VPWR
+ VPWR __dut__._1273_/X sky130_fd_sc_hd__a21o_4
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1104__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_221_ _292_/Q _220_/A _222_/A VGND VGND VPWR VPWR _295_/D sky130_fd_sc_hd__o21a_4
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_152_ _302_/Q VGND VGND VPWR VPWR _154_/C sky130_fd_sc_hd__inv_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0988_ __dut__._1378_/A __dut__._1910_/Q VGND VGND VPWR VPWR __dut__._0988_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_2_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1609_ __dut__._1543_/Y mc[24] __dut__._1608_/X VGND VGND VPWR VPWR __dut__._1609_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1059__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1_0___dut__.__uuf__.__clk_source__ clkbuf_3_1_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_4_3_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_41_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1231__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1684__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2060_ __dut__.__uuf__._2065_/CLK __dut__._1109_/X __dut__.__uuf__._1593_/X
+ VGND VGND VPWR VPWR __dut__._1110_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1844__CLK __dut__._1899_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1913_ __dut__.__uuf__._1906_/Y __dut__.__uuf__._1907_/Y __dut__.__uuf__._1906_/Y
+ __dut__.__uuf__._1907_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1914_/C sky130_fd_sc_hd__a2bb2o_4
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1844_ __dut__.__uuf__._1841_/Y __dut__.__uuf__._1842_/Y __dut__.__uuf__._1798_/X
+ __dut__.__uuf__._1848_/B VGND VGND VPWR VPWR __dut__.__uuf__._1844_/X sky130_fd_sc_hd__o22a_4
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1775_ __dut__._1044_/B VGND VGND VPWR VPWR __dut__.__uuf__._1775_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1773__A2 mp[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._0911_ __dut__._1383_/A1 prod[52] __dut__._0910_/X VGND VGND VPWR VPWR __dut__._1872_/D
+ sky130_fd_sc_hd__a21o_4
X__dut__._1891_ __dut__._1902_/CLK __dut__._1891_/D __dut__._1438_/Y VGND VGND VPWR
+ VPWR __dut__._1891_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1594__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1209_ __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR __dut__.__uuf__._1209_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._2189_ __dut__.__uuf__._2194_/CLK __dut__._1367_/X __dut__.__uuf__._1120_/X
+ VGND VGND VPWR VPWR prod[49] sky130_fd_sc_hd__dfrtp_4
XFILLER_74_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1325_ __dut__._1325_/A1 __dut__._1325_/A2 __dut__._1324_/X VGND VGND VPWR
+ VPWR __dut__._1325_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_66_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1256_ __dut__._1786_/A __dut__._1256_/B VGND VGND VPWR VPWR __dut__._1256_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__.__uuf__._2105__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_90_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1187_ __dut__._1187_/A1 __dut__._1187_/A2 __dut__._1186_/X VGND VGND VPWR
+ VPWR __dut__._1187_/X sky130_fd_sc_hd__a21o_4
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_204_ _246_/Q VGND VGND VPWR VPWR _204_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1213__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_135_ _308_/Q _231_/A VGND VGND VPWR VPWR _135_/X sky130_fd_sc_hd__and2_4
XFILLER_99_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_15_0_tck clkbuf_3_7_0_tck/X VGND VGND VPWR VPWR __dut__._1915_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA___dut__._1867__CLK __dut__._1915_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1864__A __dut__._1557_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_128_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._1560_ __dut__._1653_/X __dut__.__uuf__._1078_/A __dut__._1148_/B
+ __dut__.__uuf__._1660_/A VGND VGND VPWR VPWR __dut__.__uuf__._1560_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1491_ __dut__.__uuf__._1575_/A VGND VGND VPWR VPWR __dut__.__uuf__._1508_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_88_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2112_ __dut__.__uuf__._2114_/CLK __dut__._1213_/X __dut__.__uuf__._1409_/X
+ VGND VGND VPWR VPWR __dut__._1214_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__.__uuf__._2043_ __dut__.__uuf__._2043_/CLK __dut__._1075_/X __dut__.__uuf__._1615_/X
+ VGND VGND VPWR VPWR __dut__._1076_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1110_ __dut__._1678_/A __dut__._1110_/B VGND VGND VPWR VPWR __dut__._1110_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1041_ __dut__._1647_/A1 __dut__._1041_/A2 __dut__._1040_/X VGND VGND VPWR
+ VPWR __dut__._1041_/X sky130_fd_sc_hd__a21o_4
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1827_ __dut__.__uuf__._1826_/X __dut__.__uuf__._1825_/B __dut__.__uuf__._1825_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1828_/C sky130_fd_sc_hd__o21ai_4
X__dut__.__uuf__._1758_ __dut__.__uuf__._1868_/A VGND VGND VPWR VPWR __dut__.__uuf__._1804_/A
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1689_ __dut__.__uuf__._1683_/Y __dut__.__uuf__._1684_/Y __dut__.__uuf__._1660_/X
+ __dut__.__uuf__._1688_/X VGND VGND VPWR VPWR __dut__.__uuf__._1690_/A sky130_fd_sc_hd__a211o_4
X__dut__._1874_ __dut__._1917_/CLK __dut__._1874_/D __dut__._1455_/Y VGND VGND VPWR
+ VPWR __dut__._1874_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_3_4_0_tck clkbuf_3_5_0_tck/A VGND VGND VPWR VPWR clkbuf_4_9_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1308_ __dut__._1308_/A prod[19] VGND VGND VPWR VPWR __dut__._1308_/X sky130_fd_sc_hd__and2_4
X__dut__._1239_ __dut__._1787_/A1 __dut__._1239_/A2 __dut__._1238_/X VGND VGND VPWR
+ VPWR __dut__._1239_/X sky130_fd_sc_hd__a21o_4
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1499__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1737__A2 mp[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1673__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1612_ __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR __dut__.__uuf__._1637_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1202__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1543_ __dut__.__uuf__._1550_/A VGND VGND VPWR VPWR __dut__.__uuf__._1543_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1474_ __dut__._1745_/X __dut__.__uuf__._1472_/X __dut__._1190_/B
+ __dut__.__uuf__._1473_/X VGND VGND VPWR VPWR __dut__.__uuf__._1474_/X sky130_fd_sc_hd__o22a_4
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1590_ __dut__._1590_/A __dut__._1790_/Q VGND VGND VPWR VPWR __dut__._1590_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2026_ __dut__.__uuf__._2043_/CLK __dut__._1041_/X __dut__.__uuf__._1635_/X
+ VGND VGND VPWR VPWR __dut__._1042_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._1079__A2 __dut__.__uuf__._2003_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1024_ __dut__._1128_/A __dut__._1024_/B VGND VGND VPWR VPWR __dut__._1024_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_29_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1857_ __dut__._1883_/CLK __dut__._1857_/D __dut__._1472_/Y VGND VGND VPWR
+ VPWR __dut__._1857_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1788_ __dut__._1788_/A __dut__._1851_/Q VGND VGND VPWR VPWR __dut__._1788_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1782__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1190_ __dut__.__uuf__._1190_/A VGND VGND VPWR VPWR __dut__.__uuf__._1249_/A
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1692__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1526_ __dut__.__uuf__._1566_/A VGND VGND VPWR VPWR __dut__.__uuf__._1526_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1711_ __dut__._1719_/A1 __dut__._1709_/X __dut__._1710_/X VGND VGND VPWR
+ VPWR __dut__._1831_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1457_ __dut__.__uuf__._1443_/X __dut__.__uuf__._1437_/X __dut__._1196_/B
+ __dut__.__uuf__._1449_/X __dut__.__uuf__._1456_/X VGND VGND VPWR VPWR __dut__._1195_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__._1642_ __dut__._1642_/A __dut__._1813_/Q VGND VGND VPWR VPWR __dut__._1642_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1388_ __dut__.__uuf__._1393_/A VGND VGND VPWR VPWR __dut__.__uuf__._1388_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1573_ __dut__._1543_/Y mc[16] __dut__._1572_/X VGND VGND VPWR VPWR __dut__._1573_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1637__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2009_ __dut__.__uuf__._2114_/CLK __dut__._1007_/X __dut__.__uuf__._1655_/X
+ VGND VGND VPWR VPWR __dut__._1008_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_82_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0946__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1007_ __dut__._1787_/A1 __dut__._1007_/A2 __dut__._1006_/X VGND VGND VPWR
+ VPWR __dut__._1007_/X sky130_fd_sc_hd__a21o_4
X__dut__._1909_ __dut__._1917_/CLK __dut__._1909_/D __dut__._1420_/Y VGND VGND VPWR
+ VPWR __dut__._1909_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_psn_inst_psn_buff_110_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1311_ __dut__.__uuf__._1316_/A VGND VGND VPWR VPWR __dut__.__uuf__._1311_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1242_ __dut__.__uuf__._1466_/A VGND VGND VPWR VPWR __dut__.__uuf__._1242_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1173_ __dut__.__uuf__._1168_/X __dut__.__uuf__._1165_/X prod[31]
+ prod[32] __dut__.__uuf__._1160_/X VGND VGND VPWR VPWR __dut__._1331_/A2 sky130_fd_sc_hd__a32o_4
XANTENNA___dut__._1619__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1509_ __dut__.__uuf__._1551_/A VGND VGND VPWR VPWR __dut__.__uuf__._1509_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1625_ __dut__._1543_/Y mc[28] __dut__._1624_/X VGND VGND VPWR VPWR __dut__._1625_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_96_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1556_ __dut__._1788_/A __dut__._1793_/Q VGND VGND VPWR VPWR __dut__._1556_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1487_ rst VGND VGND VPWR VPWR __dut__._1487_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_297_ _306_/CLK _297_/D trst VGND VGND VPWR VPWR _297_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_5_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_158_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2011__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2161__CLK __dut__.__uuf__._2210_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1860_ __dut__.__uuf__._1826_/X __dut__.__uuf__._1859_/B __dut__.__uuf__._1859_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1861_/C sky130_fd_sc_hd__o21ai_4
XFILLER_17_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1791_ __dut__.__uuf__._1791_/A VGND VGND VPWR VPWR __dut__._1053_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1210__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1225_ __dut__.__uuf__._1233_/A VGND VGND VPWR VPWR __dut__.__uuf__._1225_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1156_ __dut__.__uuf__._1153_/X __dut__.__uuf__._1149_/X prod[37]
+ prod[38] __dut__.__uuf__._1145_/X VGND VGND VPWR VPWR __dut__._1343_/A2 sky130_fd_sc_hd__a32o_4
X__dut__._1410_ __dut__._1788_/A __dut__._1410_/B VGND VGND VPWR VPWR __dut__._1410_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1341_ __dut__._1341_/A1 __dut__._1341_/A2 __dut__._1340_/X VGND VGND VPWR
+ VPWR __dut__._1341_/X sky130_fd_sc_hd__a21o_4
XFILLER_47_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1087_ __dut__.__uuf__._2008_/A VGND VGND VPWR VPWR __dut__.__uuf__._1099_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_55_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1272_ __dut__._1272_/A prod[1] VGND VGND VPWR VPWR __dut__._1272_/X sky130_fd_sc_hd__and2_4
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1989_ __dut__.__uuf__._1692_/A __dut__.__uuf__._1988_/B __dut__.__uuf__._1988_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1990_/C sky130_fd_sc_hd__o21ai_4
X_220_ _220_/A _225_/B VGND VGND VPWR VPWR _294_/D sky130_fd_sc_hd__and2_4
X_151_ _312_/Q VGND VGND VPWR VPWR _238_/A sky130_fd_sc_hd__inv_2
XANTENNA_psn_inst_psn_buff_11_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1120__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0987_ __dut__._1339_/A1 prod[25] __dut__._0986_/X VGND VGND VPWR VPWR __dut__._1910_/D
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__.__uuf__._2034__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1608_ __dut__._1788_/A __dut__._1806_/Q VGND VGND VPWR VPWR __dut__._1608_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA__315__CLK _194_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1539_ rst VGND VGND VPWR VPWR __dut__._1539_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1796__CLK __dut__._1410_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1912_ __dut__.__uuf__._1912_/A VGND VGND VPWR VPWR __dut__._1097_/A2
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1843_ __dut__._1565_/X VGND VGND VPWR VPWR __dut__.__uuf__._1848_/B
+ sky130_fd_sc_hd__inv_2
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1774_ __dut__._1050_/B VGND VGND VPWR VPWR __dut__.__uuf__._1774_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._0910_ __dut__._1378_/A __dut__._1871_/Q VGND VGND VPWR VPWR __dut__._0910_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1890_ __dut__._1902_/CLK __dut__._1890_/D __dut__._1439_/Y VGND VGND VPWR
+ VPWR __dut__._1890_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1208_ __dut__.__uuf__._1218_/A VGND VGND VPWR VPWR __dut__.__uuf__._1208_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._2188_ __dut__.__uuf__._2194_/CLK __dut__._1365_/X __dut__.__uuf__._1123_/X
+ VGND VGND VPWR VPWR prod[48] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1139_ __dut__.__uuf__._1138_/X __dut__.__uuf__._1135_/X prod[43]
+ prod[44] __dut__.__uuf__._1131_/X VGND VGND VPWR VPWR __dut__._1355_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1324_ __dut__._1324_/A prod[27] VGND VGND VPWR VPWR __dut__._1324_/X sky130_fd_sc_hd__and2_4
X__dut__._1255_ __dut__._1787_/A1 __dut__._1255_/A2 __dut__._1254_/X VGND VGND VPWR
+ VPWR __dut__._1255_/X sky130_fd_sc_hd__a21o_4
XANTENNA_psn_inst_psn_buff_59_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1186_ __dut__._1770_/A __dut__._1186_/B VGND VGND VPWR VPWR __dut__._1186_/X
+ sky130_fd_sc_hd__and2_4
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._0954__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_203_ _203_/A VGND VGND VPWR VPWR _203_/X sky130_fd_sc_hd__buf_2
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_134_ _134_/A VGND VGND VPWR VPWR _313_/D sky130_fd_sc_hd__inv_2
XFILLER_99_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._0864__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1490_ __dut__.__uuf__._1612_/A VGND VGND VPWR VPWR __dut__.__uuf__._1575_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2111_ __dut__.__uuf__._2114_/CLK __dut__._1211_/X __dut__.__uuf__._1413_/X
+ VGND VGND VPWR VPWR __dut__._1212_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2042_ __dut__.__uuf__._2043_/CLK __dut__._1073_/X __dut__.__uuf__._1616_/X
+ VGND VGND VPWR VPWR __dut__._1074_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__._1040_ __dut__._1626_/A __dut__._1040_/B VGND VGND VPWR VPWR __dut__._1040_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_100_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1826_ __dut__.__uuf__._1936_/A VGND VGND VPWR VPWR __dut__.__uuf__._1826_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1757_ __dut__.__uuf__._1757_/A VGND VGND VPWR VPWR __dut__._1041_/A2
+ sky130_fd_sc_hd__inv_2
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1688_ __dut__.__uuf__._1683_/Y __dut__.__uuf__._1684_/Y __dut__.__uuf__._1686_/X
+ __dut__.__uuf__._1692_/B VGND VGND VPWR VPWR __dut__.__uuf__._1688_/X sky130_fd_sc_hd__o22a_4
X__dut__._1873_ __dut__._1917_/CLK __dut__._1873_/D __dut__._1456_/Y VGND VGND VPWR
+ VPWR __dut__._1873_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1131__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__._1307_ __dut__._1319_/A1 __dut__._1307_/A2 __dut__._1306_/X VGND VGND VPWR
+ VPWR __dut__._1307_/X sky130_fd_sc_hd__a21o_4
X__dut__._1238_ __dut__._1786_/A __dut__._1238_/B VGND VGND VPWR VPWR __dut__._1238_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_31_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1169_ __dut__._1647_/A1 __dut__._1169_/A2 __dut__._1168_/X VGND VGND VPWR
+ VPWR __dut__._1169_/X sky130_fd_sc_hd__a21o_4
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1834__CLK __dut__._1410_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1875__A __dut__._1553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1673__A2 mp[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_140_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1611_ __dut__.__uuf__._1611_/A VGND VGND VPWR VPWR __dut__.__uuf__._1611_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1542_ __dut__.__uuf__._1530_/X __dut__.__uuf__._1526_/X __dut__._1156_/B
+ __dut__.__uuf__._1535_/X __dut__.__uuf__._1541_/X VGND VGND VPWR VPWR __dut__._1155_/A2
+ sky130_fd_sc_hd__a32o_4
XANTENNA___dut__.__uuf__._1260__A3 prod[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1473_ __dut__.__uuf__._1495_/A VGND VGND VPWR VPWR __dut__.__uuf__._1473_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_89_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1361__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2025_ __dut__.__uuf__._2043_/CLK __dut__._1039_/X __dut__.__uuf__._1636_/X
+ VGND VGND VPWR VPWR __dut__._1040_/B sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__._1113__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__.__uuf__._1079__A3 prod[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_14_0_tck clkbuf_3_7_0_tck/X VGND VGND VPWR VPWR __dut__._1917_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_25_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__._1023_ __dut__._1129_/A1 __dut__._1023_/A2 __dut__._1022_/X VGND VGND VPWR
+ VPWR __dut__._1023_/X sky130_fd_sc_hd__a21o_4
XFILLER_25_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X__dut__.__uuf__._1809_ __dut__._1577_/X VGND VGND VPWR VPWR __dut__.__uuf__._1815_/B
+ sky130_fd_sc_hd__inv_2
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1856_ __dut__._1919_/CLK __dut__._1856_/D __dut__._1473_/Y VGND VGND VPWR
+ VPWR __dut__._1856_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1787_ __dut__._1787_/A1 __dut__._1785_/X __dut__._1786_/X VGND VGND VPWR
+ VPWR __dut__._1850_/D sky130_fd_sc_hd__a21o_4
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1591__A1 __dut__._1647_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2118__CLK __dut__.__uuf__._2119_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_98_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3_0_tck clkbuf_3_3_0_tck/A VGND VGND VPWR VPWR clkbuf_4_7_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0909__A1 __dut__._1383_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1525_ __dut__.__uuf__._1529_/A VGND VGND VPWR VPWR __dut__.__uuf__._1525_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1710_ __dut__._1766_/A __dut__._1830_/Q VGND VGND VPWR VPWR __dut__._1710_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1456_ __dut__._1761_/X __dut__.__uuf__._1451_/X __dut__._1198_/B
+ __dut__.__uuf__._1452_/X VGND VGND VPWR VPWR __dut__.__uuf__._1456_/X sky130_fd_sc_hd__o22a_4
X__dut__._1641_ __dut__._1543_/Y mc[31] __dut__._1640_/X VGND VGND VPWR VPWR __dut__._1641_/X
+ sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1387_ __dut__.__uuf__._1380_/X __dut__.__uuf__._1386_/X __dut__._1224_/B
+ __dut__.__uuf__._1380_/X VGND VGND VPWR VPWR __dut__._1223_/A2 sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1572_ __dut__._1788_/A __dut__._1797_/Q VGND VGND VPWR VPWR __dut__._1572_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2008_ __dut__.__uuf__._2008_/A VGND VGND VPWR VPWR __dut__.__uuf__._2008_/X
+ sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1637__A2 mc[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_41_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X__dut__._1006_ __dut__._1786_/A __dut__._1850_/Q VGND VGND VPWR VPWR __dut__._1006_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._1573__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1908_ __dut__._1919_/CLK __dut__._1908_/D __dut__._1421_/Y VGND VGND VPWR
+ VPWR __dut__._1908_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1839_ __dut__._1899_/CLK __dut__._1839_/D __dut__._1490_/Y VGND VGND VPWR
+ VPWR __dut__._1839_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0872__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_103_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1310_ __dut__.__uuf__._1303_/X __dut__.__uuf__._1309_/X __dut__._1254_/B
+ __dut__.__uuf__._1303_/X VGND VGND VPWR VPWR __dut__._1253_/A2 sky130_fd_sc_hd__a2bb2o_4
X__dut__.__uuf__._1241_ __dut__.__uuf__._1248_/A VGND VGND VPWR VPWR __dut__.__uuf__._1241_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1172_ __dut__.__uuf__._1174_/A VGND VGND VPWR VPWR __dut__.__uuf__._1172_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1208__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1619__A2 __dut__._1617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA___dut__._1555__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1508_ __dut__.__uuf__._1508_/A VGND VGND VPWR VPWR __dut__.__uuf__._1508_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1439_ __dut__.__uuf__._1536_/A VGND VGND VPWR VPWR __dut__.__uuf__._1946_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1624_ __dut__._1788_/A __dut__._1810_/Q VGND VGND VPWR VPWR __dut__._1624_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA_psn_inst_psn_buff_89_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1555_ __dut__._1767_/A1 __dut__._1553_/X __dut__._1554_/X VGND VGND VPWR
+ VPWR __dut__._1792_/D sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1118__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1486_ rst VGND VGND VPWR VPWR __dut__._1486_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1788__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_296_ _313_/CLK _296_/D trst VGND VGND VPWR VPWR _296_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1790_ __dut__.__uuf__._1786_/Y __dut__.__uuf__._1787_/Y __dut__.__uuf__._1776_/X
+ __dut__.__uuf__._1789_/X VGND VGND VPWR VPWR __dut__.__uuf__._1791_/A sky130_fd_sc_hd__a211o_4
XFILLER_20_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1698__A __dut__._1766_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1785__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1918__CLK __dut__._1919_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1224_ __dut__.__uuf__._1212_/X __dut__.__uuf__._1223_/X prod[14]
+ prod[15] __dut__.__uuf__._1219_/X VGND VGND VPWR VPWR __dut__._1297_/A2 sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1155_ __dut__.__uuf__._1159_/A VGND VGND VPWR VPWR __dut__.__uuf__._1155_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1086_ __dut__.__uuf__._1075_/X __dut__.__uuf__._2003_/A prod[60]
+ prod[61] __dut__.__uuf__._1085_/X VGND VGND VPWR VPWR __dut__._1389_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_86_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1340_ __dut__._1340_/A prod[35] VGND VGND VPWR VPWR __dut__._1340_/X sky130_fd_sc_hd__and2_4
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1271_ __dut__._1273_/A1 __dut__._1271_/A2 __dut__._1270_/X VGND VGND VPWR
+ VPWR __dut__._1271_/X sky130_fd_sc_hd__a21o_4
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1988_ __dut__.__uuf__._2001_/A __dut__.__uuf__._1988_/B __dut__.__uuf__._1988_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1990_/B sky130_fd_sc_hd__or3_4
X_150_ _146_/Y _296_/Q _308_/Q _307_/Q _220_/A VGND VGND VPWR VPWR _307_/D sky130_fd_sc_hd__o32a_4
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0986_ __dut__._1378_/A __dut__._1909_/Q VGND VGND VPWR VPWR __dut__._0986_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_2_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1607_ __dut__._1767_/A1 __dut__._1605_/X __dut__._1606_/X VGND VGND VPWR
+ VPWR __dut__._1805_/D sky130_fd_sc_hd__a21o_4
X__dut__._1538_ rst VGND VGND VPWR VPWR __dut__._1538_/Y sky130_fd_sc_hd__inv_2
X__dut__._1469_ rst VGND VGND VPWR VPWR __dut__._1469_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1767__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_279_ _314_/CLK _279_/D VGND VGND VPWR VPWR _279_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_170_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1911_ __dut__.__uuf__._1906_/Y __dut__.__uuf__._1907_/Y __dut__.__uuf__._1886_/X
+ __dut__.__uuf__._1910_/X VGND VGND VPWR VPWR __dut__.__uuf__._1912_/A sky130_fd_sc_hd__a211o_4
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1842_ __dut__._1068_/B VGND VGND VPWR VPWR __dut__.__uuf__._1842_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1773_ __dut__.__uuf__._1773_/A __dut__.__uuf__._1773_/B __dut__.__uuf__._1773_/C
+ VGND VGND VPWR VPWR __dut__._1043_/A2 sky130_fd_sc_hd__and3_4
XANTENNA___dut__._1890__CLK __dut__._1902_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0___dut__.__uuf__.__clk_source__ clkbuf_2_3_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0___dut__.__uuf__.__clk_source__/A sky130_fd_sc_hd__clkbuf_1
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2187_ __dut__.__uuf__._2194_/CLK __dut__._1363_/X __dut__.__uuf__._1126_/X
+ VGND VGND VPWR VPWR prod[47] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1207_ __dut__.__uuf__._1236_/A VGND VGND VPWR VPWR __dut__.__uuf__._1218_/A
+ sky130_fd_sc_hd__buf_2
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__.__uuf__._1138_ __dut__.__uuf__._1138_/A VGND VGND VPWR VPWR __dut__.__uuf__._1138_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1323_ __dut__._1323_/A1 __dut__._1323_/A2 __dut__._1322_/X VGND VGND VPWR
+ VPWR __dut__._1323_/X sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1069_ __dut__.__uuf__._1190_/A VGND VGND VPWR VPWR __dut__.__uuf__._1069_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1254_ __dut__._1786_/A __dut__._1254_/B VGND VGND VPWR VPWR __dut__._1254_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_70_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1185_ __dut__._1187_/A1 __dut__._1185_/A2 __dut__._1184_/X VGND VGND VPWR
+ VPWR __dut__._1185_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1749__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_202_ _203_/A VGND VGND VPWR VPWR _202_/X sky130_fd_sc_hd__buf_2
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_133_ _131_/Y _231_/A _132_/Y _128_/X VGND VGND VPWR VPWR _134_/A sky130_fd_sc_hd__a211o_4
X__dut__._0969_ __dut__._1319_/A1 prod[16] __dut__._0968_/X VGND VGND VPWR VPWR __dut__._1901_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_78_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2110_ __dut__.__uuf__._2138_/CLK __dut__._1209_/X __dut__.__uuf__._1418_/X
+ VGND VGND VPWR VPWR __dut__._1210_/B sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._2041_ __dut__.__uuf__._2043_/CLK __dut__._1071_/X __dut__.__uuf__._1617_/X
+ VGND VGND VPWR VPWR __dut__._1072_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1216__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1825_ __dut__.__uuf__._1859_/A __dut__.__uuf__._1825_/B __dut__.__uuf__._1825_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1828_/B sky130_fd_sc_hd__or3_4
XFILLER_100_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1756_ __dut__.__uuf__._1752_/Y __dut__.__uuf__._1753_/Y __dut__.__uuf__._1721_/X
+ __dut__.__uuf__._1755_/X VGND VGND VPWR VPWR __dut__.__uuf__._1757_/A sky130_fd_sc_hd__a211o_4
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1687_ __dut__._1625_/X VGND VGND VPWR VPWR __dut__.__uuf__._1692_/B
+ sky130_fd_sc_hd__inv_2
X__dut__._1872_ __dut__._1915_/CLK __dut__._1872_/D __dut__._1457_/Y VGND VGND VPWR
+ VPWR __dut__._1872_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_48_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_71_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1126__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1306_ __dut__._1308_/A prod[18] VGND VGND VPWR VPWR __dut__._1306_/X sky130_fd_sc_hd__and2_4
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1237_ __dut__._1787_/A1 __dut__._1237_/A2 __dut__._1236_/X VGND VGND VPWR
+ VPWR __dut__._1237_/X sky130_fd_sc_hd__a21o_4
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1168_ __dut__._1174_/A __dut__._1168_/B VGND VGND VPWR VPWR __dut__._1168_/X
+ sky130_fd_sc_hd__and2_4
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1099_ __dut__._1129_/A1 __dut__._1099_/A2 __dut__._1098_/X VGND VGND VPWR
+ VPWR __dut__._1099_/X sky130_fd_sc_hd__a21o_4
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1036__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1891__A __dut__.__uuf__._1946_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2047__CLK __dut__.__uuf__._2049_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_psn_inst_psn_buff_133_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1610_ __dut__.__uuf__._1611_/A VGND VGND VPWR VPWR __dut__.__uuf__._1610_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1541_ __dut__._1673_/X __dut__.__uuf__._1536_/X __dut__._1158_/B
+ __dut__.__uuf__._1537_/X VGND VGND VPWR VPWR __dut__.__uuf__._1541_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1472_ __dut__.__uuf__._1536_/A VGND VGND VPWR VPWR __dut__.__uuf__._1472_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2024_ __dut__.__uuf__._2043_/CLK __dut__._1037_/X __dut__.__uuf__._1638_/X
+ VGND VGND VPWR VPWR __dut__._1038_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_57_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1022_ __dut__._1128_/A __dut__._1022_/B VGND VGND VPWR VPWR __dut__._1022_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_71_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X__dut__.__uuf__._1808_ __dut__._1056_/B VGND VGND VPWR VPWR __dut__.__uuf__._1808_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._0927__A2 prod[60] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1739_ __dut__.__uuf__._1715_/X __dut__.__uuf__._1738_/B __dut__.__uuf__._1738_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1740_/C sky130_fd_sc_hd__o21ai_4
X__dut__._1855_ __dut__._1919_/CLK __dut__._1855_/D __dut__._1474_/Y VGND VGND VPWR
+ VPWR __dut__._1855_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1786_ __dut__._1786_/A __dut__._1849_/Q VGND VGND VPWR VPWR __dut__._1786_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_96_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_5_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0863__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1031__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1524_ __dut__.__uuf__._1509_/X __dut__.__uuf__._1505_/X __dut__._1164_/B
+ __dut__.__uuf__._1514_/X __dut__.__uuf__._1523_/X VGND VGND VPWR VPWR __dut__._1163_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1455_ __dut__.__uuf__._1465_/A VGND VGND VPWR VPWR __dut__.__uuf__._1455_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1640_ __dut__._1788_/A __dut__._1814_/Q VGND VGND VPWR VPWR __dut__._1640_/X
+ sky130_fd_sc_hd__and2_4
X__dut__.__uuf__._1386_ __dut__.__uuf__._1385_/Y __dut__.__uuf__._1375_/X __dut__.__uuf__._1376_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1386_/X sky130_fd_sc_hd__o21a_4
XFILLER_89_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1571_ __dut__._1767_/A1 __dut__._1569_/X __dut__._1570_/X VGND VGND VPWR
+ VPWR __dut__._1796_/D sky130_fd_sc_hd__a21o_4
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2007_ done __dut__.__uuf__._2006_/Y __dut__._1785_/X VGND VGND VPWR
+ VPWR __dut__._1137_/A2 sky130_fd_sc_hd__o21a_4
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_34_A psn_inst_psn_buff_49/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1005_ __dut__._1005_/A1 prod[34] __dut__._1004_/X VGND VGND VPWR VPWR __dut__._1919_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1573__A2 mc[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1907_ __dut__._1919_/CLK __dut__._1907_/D __dut__._1422_/Y VGND VGND VPWR
+ VPWR __dut__._1907_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1838_ __dut__._1899_/CLK __dut__._1838_/D __dut__._1491_/Y VGND VGND VPWR
+ VPWR __dut__._1838_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1769_ __dut__._1543_/Y mp[28] __dut__._1768_/X VGND VGND VPWR VPWR __dut__._1769_/X
+ sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1089__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1261__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1013__A1 __dut__._1129_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_4_0___dut__.__uuf__.__clk_source__ clkbuf_4_5_0___dut__.__uuf__.__clk_source__/A
+ VGND VGND VPWR VPWR __dut__.__uuf__._2043_/CLK sky130_fd_sc_hd__clkbuf_1
X__dut__.__uuf__._1240_ __dut__.__uuf__._1227_/X __dut__.__uuf__._1239_/X prod[9]
+ prod[10] __dut__.__uuf__._1234_/X VGND VGND VPWR VPWR __dut__._1287_/A2 sky130_fd_sc_hd__a32o_4
Xclkbuf_4_13_0_tck clkbuf_3_6_0_tck/X VGND VGND VPWR VPWR __dut__._1899_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1171_ __dut__.__uuf__._1168_/X __dut__.__uuf__._1165_/X prod[32]
+ prod[33] __dut__.__uuf__._1160_/X VGND VGND VPWR VPWR __dut__._1333_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_101_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1224__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA___dut__._1555__A2 __dut__._1553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1507_ __dut__.__uuf__._1487_/X __dut__.__uuf__._1505_/X __dut__._1172_/B
+ __dut__.__uuf__._1493_/X __dut__.__uuf__._1506_/X VGND VGND VPWR VPWR __dut__._1171_/A2
+ sky130_fd_sc_hd__a32o_4
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1438_ __dut__.__uuf__._1438_/A VGND VGND VPWR VPWR __dut__.__uuf__._1536_/A
+ sky130_fd_sc_hd__buf_2
X__dut__._1623_ __dut__._1767_/A1 __dut__._1621_/X __dut__._1622_/X VGND VGND VPWR
+ VPWR __dut__._1809_/D sky130_fd_sc_hd__a21o_4
X__dut__.__uuf__._1369_ __dut__.__uuf__._1368_/Y __dut__.__uuf__._1349_/X __dut__.__uuf__._1350_/X
+ VGND VGND VPWR VPWR __dut__.__uuf__._1369_/X sky130_fd_sc_hd__o21a_4
X__dut__._1554_ __dut__._1766_/A __dut__._1791_/Q VGND VGND VPWR VPWR __dut__._1554_/X
+ sky130_fd_sc_hd__and2_4
X__dut__._1485_ rst VGND VGND VPWR VPWR __dut__._1485_/Y sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1134__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2108__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1243__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_295_ _314_/CLK _295_/D trst VGND VGND VPWR VPWR _295_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_tck clkbuf_3_3_0_tck/A VGND VGND VPWR VPWR clkbuf_4_5_0_tck/A sky130_fd_sc_hd__clkbuf_1
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1785__A2 start VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X__dut__.__uuf__._1223_ __dut__.__uuf__._1223_/A VGND VGND VPWR VPWR __dut__.__uuf__._1223_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_101_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1154_ __dut__.__uuf__._1153_/X __dut__.__uuf__._1149_/X prod[38]
+ prod[39] __dut__.__uuf__._1145_/X VGND VGND VPWR VPWR __dut__._1345_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_59_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1085_ __dut__.__uuf__._1100_/A VGND VGND VPWR VPWR __dut__.__uuf__._1085_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1270_ __dut__._1270_/A prod[0] VGND VGND VPWR VPWR __dut__._1270_/X sky130_fd_sc_hd__and2_4
XFILLER_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__300__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__.__uuf__._1987_ __dut__.__uuf__._1981_/Y __dut__.__uuf__._1982_/Y __dut__.__uuf__._1981_/Y
+ __dut__.__uuf__._1982_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1988_/C sky130_fd_sc_hd__a2bb2o_4
XANTENNA___dut__._1225__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0985_ __dut__._1339_/A1 prod[24] __dut__._0984_/X VGND VGND VPWR VPWR __dut__._1909_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1606_ __dut__._1766_/A __dut__._1804_/Q VGND VGND VPWR VPWR __dut__._1606_/X
+ sky130_fd_sc_hd__and2_4
XANTENNA___dut__._0968__A __dut__._1770_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1537_ rst VGND VGND VPWR VPWR __dut__._1537_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1468_ rst VGND VGND VPWR VPWR __dut__._1468_/Y sky130_fd_sc_hd__inv_2
X__dut__._1399_ __dut__._1787_/A1 __dut__._1399_/A2 __dut__._1398_/X VGND VGND VPWR
+ VPWR __dut__._1399_/X sky130_fd_sc_hd__a21o_4
XANTENNA___dut__._1767__A2 __dut__._1765_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_278_ _314_/CLK _278_/D VGND VGND VPWR VPWR _278_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_163_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1910_ __dut__.__uuf__._1906_/Y __dut__.__uuf__._1907_/Y __dut__.__uuf__._1908_/X
+ __dut__.__uuf__._1914_/B VGND VGND VPWR VPWR __dut__.__uuf__._1910_/X sky130_fd_sc_hd__o22a_4
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1841_ __dut__._1074_/B VGND VGND VPWR VPWR __dut__.__uuf__._1841_/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA___dut__._1207__A1 __dut__._1787_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1502__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1772_ __dut__.__uuf__._1771_/X __dut__.__uuf__._1770_/B __dut__.__uuf__._1770_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1773_/C sky130_fd_sc_hd__o21ai_4
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2186_ __dut__.__uuf__._2194_/CLK __dut__._1361_/X __dut__.__uuf__._1128_/X
+ VGND VGND VPWR VPWR prod[46] sky130_fd_sc_hd__dfrtp_4
X__dut__.__uuf__._1206_ __dut__.__uuf__._1198_/X __dut__.__uuf__._1195_/X prod[20]
+ prod[21] __dut__.__uuf__._1205_/X VGND VGND VPWR VPWR __dut__._1309_/A2 sky130_fd_sc_hd__a32o_4
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1137_ __dut__.__uuf__._1144_/A VGND VGND VPWR VPWR __dut__.__uuf__._1137_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_74_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1068_ __dut__.__uuf__._1084_/A VGND VGND VPWR VPWR __dut__.__uuf__._1068_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1322_ __dut__._1324_/A prod[26] VGND VGND VPWR VPWR __dut__._1322_/X sky130_fd_sc_hd__and2_4
X__dut__._1253_ __dut__._1787_/A1 __dut__._1253_/A2 __dut__._1252_/X VGND VGND VPWR
+ VPWR __dut__._1253_/X sky130_fd_sc_hd__a21o_4
XFILLER_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1412__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1184_ __dut__._1770_/A __dut__._1184_/B VGND VGND VPWR VPWR __dut__._1184_/X
+ sky130_fd_sc_hd__and2_4
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_201_ _203_/A VGND VGND VPWR VPWR _201_/X sky130_fd_sc_hd__buf_2
XANTENNA___dut__._1749__A2 mp[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_132_ _313_/Q _231_/A VGND VGND VPWR VPWR _132_/Y sky130_fd_sc_hd__nor2_4
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0968_ __dut__._1770_/A __dut__._1900_/Q VGND VGND VPWR VPWR __dut__._0968_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._0899_ __dut__._1383_/A1 prod[46] __dut__._0898_/X VGND VGND VPWR VPWR __dut__._1866_/D
+ sky130_fd_sc_hd__a21o_4
XFILLER_78_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__293__RESET_B trst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1908__CLK __dut__._1919_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1685__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2040_ __dut__.__uuf__._2043_/CLK __dut__._1069_/X __dut__.__uuf__._1618_/X
+ VGND VGND VPWR VPWR __dut__._1070_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_96_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1232__A __dut__._1786_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1824_ __dut__.__uuf__._1818_/Y __dut__.__uuf__._1819_/Y __dut__.__uuf__._1818_/Y
+ __dut__.__uuf__._1819_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1825_/C sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1755_ __dut__.__uuf__._1752_/Y __dut__.__uuf__._1753_/Y __dut__.__uuf__._1743_/X
+ __dut__.__uuf__._1760_/B VGND VGND VPWR VPWR __dut__.__uuf__._1755_/X sky130_fd_sc_hd__o22a_4
XFILLER_20_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1686_ __dut__.__uuf__._1923_/A VGND VGND VPWR VPWR __dut__.__uuf__._1686_/X
+ sky130_fd_sc_hd__buf_2
X__dut__._1871_ __dut__._1915_/CLK __dut__._1871_/D __dut__._1458_/Y VGND VGND VPWR
+ VPWR __dut__._1871_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__._1667__A1 __dut__._1767_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2169_ __dut__.__uuf__._2169_/CLK __dut__._1327_/X __dut__.__uuf__._1179_/X
+ VGND VGND VPWR VPWR prod[29] sky130_fd_sc_hd__dfrtp_4
XFILLER_28_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_64_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__._1305_ __dut__._1319_/A1 __dut__._1305_/A2 __dut__._1304_/X VGND VGND VPWR
+ VPWR __dut__._1305_/X sky130_fd_sc_hd__a21o_4
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1236_ __dut__._1786_/A __dut__._1236_/B VGND VGND VPWR VPWR __dut__._1236_/X
+ sky130_fd_sc_hd__and2_4
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1167_ __dut__._1167_/A1 __dut__._1167_/A2 __dut__._1166_/X VGND VGND VPWR
+ VPWR __dut__._1167_/X sky130_fd_sc_hd__a21o_4
XFILLER_43_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X__dut__._1098_ __dut__._1098_/A __dut__._1098_/B VGND VGND VPWR VPWR __dut__._1098_/X
+ sky130_fd_sc_hd__and2_4
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_psn_inst_psn_buff_126_A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__._1052__A __dut__._1678_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1540_ __dut__.__uuf__._1550_/A VGND VGND VPWR VPWR __dut__.__uuf__._1540_/X
+ sky130_fd_sc_hd__buf_2
X__dut__.__uuf__._1471_ __dut__.__uuf__._1535_/A VGND VGND VPWR VPWR __dut__.__uuf__._1471_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA___dut__._1649__A1 __dut__._1543_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._2023_ __dut__.__uuf__._2049_/CLK __dut__._1035_/X __dut__.__uuf__._1639_/X
+ VGND VGND VPWR VPWR __dut__._1036_/B sky130_fd_sc_hd__dfrtp_4
XFILLER_84_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1021_ __dut__._1129_/A1 __dut__._1021_/A2 __dut__._1020_/X VGND VGND VPWR
+ VPWR __dut__._1021_/X sky130_fd_sc_hd__a21o_4
XFILLER_40_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA___dut__.__uuf__._2141__CLK __dut__.__uuf__._2208_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__.__uuf__._1807_ __dut__._1062_/B VGND VGND VPWR VPWR __dut__.__uuf__._1807_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__.__uuf__._1738_ __dut__.__uuf__._1749_/A __dut__.__uuf__._1738_/B __dut__.__uuf__._1738_/C
+ VGND VGND VPWR VPWR __dut__.__uuf__._1740_/B sky130_fd_sc_hd__or3_4
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1669_ __dut__.__uuf__._1658_/Y __dut__.__uuf__._1659_/Y __dut__.__uuf__._1658_/Y
+ __dut__.__uuf__._1659_/Y VGND VGND VPWR VPWR __dut__.__uuf__._1670_/C sky130_fd_sc_hd__a2bb2o_4
X__dut__._1854_ clkbuf_4_5_0_tck/X __dut__._1854_/D __dut__._1475_/Y VGND VGND VPWR
+ VPWR __dut__._1854_/Q sky130_fd_sc_hd__dfrtp_4
X__dut__._1785_ __dut__._1543_/Y start __dut__._1784_/X VGND VGND VPWR VPWR __dut__._1785_/X
+ sky130_fd_sc_hd__a21o_4
XFILLER_96_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0863__A2 __dut__._1789_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1219_ __dut__._1787_/A1 __dut__._1219_/A2 __dut__._1218_/X VGND VGND VPWR
+ VPWR __dut__._1219_/X sky130_fd_sc_hd__a21o_4
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA___dut__._1600__A __dut__._1788_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__.__uuf__._2014__CLK __dut__.__uuf__._2114_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._0886__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._2164__CLK __dut__.__uuf__._2164_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_66_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1510__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__.__uuf__._1523_ __dut__._1693_/X __dut__.__uuf__._1515_/X __dut__._1166_/B
+ __dut__.__uuf__._1516_/X VGND VGND VPWR VPWR __dut__.__uuf__._1523_/X sky130_fd_sc_hd__o22a_4
X__dut__.__uuf__._1454_ __dut__.__uuf__._1443_/X __dut__.__uuf__._1437_/X __dut__._1198_/B
+ __dut__.__uuf__._1449_/X __dut__.__uuf__._1453_/X VGND VGND VPWR VPWR __dut__._1197_/A2
+ sky130_fd_sc_hd__a32o_4
X__dut__.__uuf__._1385_ __dut__._1226_/B VGND VGND VPWR VPWR __dut__.__uuf__._1385_/Y
+ sky130_fd_sc_hd__inv_2
X__dut__._1570_ __dut__._1766_/A __dut__._1795_/Q VGND VGND VPWR VPWR __dut__._1570_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._2006_ __dut__.__uuf__._2006_/A VGND VGND VPWR VPWR __dut__.__uuf__._2006_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1004_ __dut__._1004_/A __dut__._1918_/Q VGND VGND VPWR VPWR __dut__._1004_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1420__A rst VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_psn_inst_psn_buff_27_A psn_inst_psn_buff_9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__._1906_ __dut__._1919_/CLK __dut__._1906_/D __dut__._1423_/Y VGND VGND VPWR
+ VPWR __dut__._1906_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA___dut__.__uuf__._2037__CLK __dut__.__uuf__._2083_/CLK VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X__dut__._1837_ __dut__._1902_/CLK __dut__._1837_/D __dut__._1492_/Y VGND VGND VPWR
+ VPWR __dut__._1837_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X__dut__._1768_ __dut__._1788_/A __dut__._1846_/Q VGND VGND VPWR VPWR __dut__._1768_/X
+ sky130_fd_sc_hd__and2_4
XFILLER_76_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X__dut__._1699_ __dut__._1719_/A1 __dut__._1697_/X __dut__._1698_/X VGND VGND VPWR
+ VPWR __dut__._1828_/D sky130_fd_sc_hd__a21o_4
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA___dut__._1799__CLK __dut__._1410_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA___dut__._1330__A __dut__._1378_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA___dut__.__uuf__._1081__B1 prod[63] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X__dut__.__uuf__._1170_ __dut__.__uuf__._1174_/A VGND VGND VPWR VPWR __dut__.__uuf__._1170_/X
+ sky130_fd_sc_hd__buf_2
XFILLER_100_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

