VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_top
  CLASS BLOCK ;
  FOREIGN user_proj_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 450.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END done
  PIN mc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END mc[0]
  PIN mc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END mc[10]
  PIN mc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END mc[11]
  PIN mc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END mc[12]
  PIN mc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END mc[13]
  PIN mc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END mc[14]
  PIN mc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END mc[15]
  PIN mc[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END mc[16]
  PIN mc[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END mc[17]
  PIN mc[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END mc[18]
  PIN mc[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END mc[19]
  PIN mc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END mc[1]
  PIN mc[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END mc[20]
  PIN mc[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END mc[21]
  PIN mc[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END mc[22]
  PIN mc[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END mc[23]
  PIN mc[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END mc[24]
  PIN mc[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END mc[25]
  PIN mc[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END mc[26]
  PIN mc[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END mc[27]
  PIN mc[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END mc[28]
  PIN mc[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END mc[29]
  PIN mc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END mc[2]
  PIN mc[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END mc[30]
  PIN mc[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END mc[31]
  PIN mc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END mc[3]
  PIN mc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END mc[4]
  PIN mc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END mc[5]
  PIN mc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END mc[6]
  PIN mc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END mc[7]
  PIN mc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END mc[8]
  PIN mc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END mc[9]
  PIN mp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END mp[0]
  PIN mp[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END mp[10]
  PIN mp[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END mp[11]
  PIN mp[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END mp[12]
  PIN mp[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END mp[13]
  PIN mp[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END mp[14]
  PIN mp[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END mp[15]
  PIN mp[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END mp[16]
  PIN mp[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END mp[17]
  PIN mp[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END mp[18]
  PIN mp[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END mp[19]
  PIN mp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END mp[1]
  PIN mp[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END mp[20]
  PIN mp[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END mp[21]
  PIN mp[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END mp[22]
  PIN mp[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END mp[23]
  PIN mp[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END mp[24]
  PIN mp[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END mp[25]
  PIN mp[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END mp[26]
  PIN mp[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END mp[27]
  PIN mp[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END mp[28]
  PIN mp[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END mp[29]
  PIN mp[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END mp[2]
  PIN mp[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END mp[30]
  PIN mp[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END mp[31]
  PIN mp[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END mp[3]
  PIN mp[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END mp[4]
  PIN mp[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END mp[5]
  PIN mp[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END mp[6]
  PIN mp[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END mp[7]
  PIN mp[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END mp[8]
  PIN mp[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END mp[9]
  PIN prod[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END prod[0]
  PIN prod[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END prod[10]
  PIN prod[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END prod[11]
  PIN prod[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END prod[12]
  PIN prod[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END prod[13]
  PIN prod[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END prod[14]
  PIN prod[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END prod[15]
  PIN prod[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END prod[16]
  PIN prod[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END prod[17]
  PIN prod[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END prod[18]
  PIN prod[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END prod[19]
  PIN prod[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END prod[1]
  PIN prod[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END prod[20]
  PIN prod[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END prod[21]
  PIN prod[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END prod[22]
  PIN prod[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END prod[23]
  PIN prod[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END prod[24]
  PIN prod[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END prod[25]
  PIN prod[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END prod[26]
  PIN prod[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END prod[27]
  PIN prod[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END prod[28]
  PIN prod[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END prod[29]
  PIN prod[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END prod[2]
  PIN prod[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END prod[30]
  PIN prod[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END prod[31]
  PIN prod[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END prod[3]
  PIN prod[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END prod[4]
  PIN prod[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END prod[5]
  PIN prod[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END prod[6]
  PIN prod[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END prod[7]
  PIN prod[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END prod[8]
  PIN prod[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END prod[9]
  PIN prod_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END prod_sel
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END rst
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END start
  PIN tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 6.840 400.000 7.440 ;
    END
  END tck
  PIN tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 88.440 400.000 89.040 ;
    END
  END tdi
  PIN tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.040 400.000 170.640 ;
    END
  END tdo
  PIN tdo_paden_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 183.640 400.000 184.240 ;
    END
  END tdo_paden_o
  PIN tie[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END tie[0]
  PIN tie[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 197.240 400.000 197.840 ;
    END
  END tie[100]
  PIN tie[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 210.840 400.000 211.440 ;
    END
  END tie[101]
  PIN tie[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 224.440 400.000 225.040 ;
    END
  END tie[102]
  PIN tie[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.720 400.000 239.320 ;
    END
  END tie[103]
  PIN tie[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 252.320 400.000 252.920 ;
    END
  END tie[104]
  PIN tie[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 265.920 400.000 266.520 ;
    END
  END tie[105]
  PIN tie[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 279.520 400.000 280.120 ;
    END
  END tie[106]
  PIN tie[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 293.120 400.000 293.720 ;
    END
  END tie[107]
  PIN tie[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.720 400.000 307.320 ;
    END
  END tie[108]
  PIN tie[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 320.320 400.000 320.920 ;
    END
  END tie[109]
  PIN tie[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END tie[10]
  PIN tie[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 446.000 11.410 450.000 ;
    END
  END tie[110]
  PIN tie[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 446.000 33.490 450.000 ;
    END
  END tie[111]
  PIN tie[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 446.000 55.570 450.000 ;
    END
  END tie[112]
  PIN tie[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 446.000 78.110 450.000 ;
    END
  END tie[113]
  PIN tie[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 446.000 100.190 450.000 ;
    END
  END tie[114]
  PIN tie[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 446.000 122.270 450.000 ;
    END
  END tie[115]
  PIN tie[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 446.000 144.810 450.000 ;
    END
  END tie[116]
  PIN tie[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 446.000 166.890 450.000 ;
    END
  END tie[117]
  PIN tie[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 446.000 188.970 450.000 ;
    END
  END tie[118]
  PIN tie[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END tie[119]
  PIN tie[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END tie[11]
  PIN tie[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END tie[120]
  PIN tie[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END tie[121]
  PIN tie[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END tie[122]
  PIN tie[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END tie[123]
  PIN tie[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END tie[124]
  PIN tie[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END tie[125]
  PIN tie[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END tie[126]
  PIN tie[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END tie[127]
  PIN tie[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END tie[128]
  PIN tie[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END tie[129]
  PIN tie[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END tie[12]
  PIN tie[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END tie[130]
  PIN tie[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END tie[131]
  PIN tie[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END tie[132]
  PIN tie[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 34.040 400.000 34.640 ;
    END
  END tie[133]
  PIN tie[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 74.840 400.000 75.440 ;
    END
  END tie[134]
  PIN tie[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 115.640 400.000 116.240 ;
    END
  END tie[135]
  PIN tie[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 156.440 400.000 157.040 ;
    END
  END tie[136]
  PIN tie[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 333.920 400.000 334.520 ;
    END
  END tie[137]
  PIN tie[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 347.520 400.000 348.120 ;
    END
  END tie[138]
  PIN tie[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 361.120 400.000 361.720 ;
    END
  END tie[139]
  PIN tie[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END tie[13]
  PIN tie[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 374.720 400.000 375.320 ;
    END
  END tie[140]
  PIN tie[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 388.320 400.000 388.920 ;
    END
  END tie[141]
  PIN tie[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 401.920 400.000 402.520 ;
    END
  END tie[142]
  PIN tie[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 415.520 400.000 416.120 ;
    END
  END tie[143]
  PIN tie[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 429.120 400.000 429.720 ;
    END
  END tie[144]
  PIN tie[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 442.720 400.000 443.320 ;
    END
  END tie[145]
  PIN tie[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 446.000 211.510 450.000 ;
    END
  END tie[146]
  PIN tie[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 446.000 233.590 450.000 ;
    END
  END tie[147]
  PIN tie[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 446.000 255.670 450.000 ;
    END
  END tie[148]
  PIN tie[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 446.000 278.210 450.000 ;
    END
  END tie[149]
  PIN tie[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END tie[14]
  PIN tie[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 446.000 300.290 450.000 ;
    END
  END tie[150]
  PIN tie[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 446.000 322.370 450.000 ;
    END
  END tie[151]
  PIN tie[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 446.000 344.910 450.000 ;
    END
  END tie[152]
  PIN tie[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 446.000 366.990 450.000 ;
    END
  END tie[153]
  PIN tie[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 446.000 389.070 450.000 ;
    END
  END tie[154]
  PIN tie[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END tie[155]
  PIN tie[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END tie[156]
  PIN tie[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END tie[157]
  PIN tie[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END tie[158]
  PIN tie[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END tie[159]
  PIN tie[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END tie[15]
  PIN tie[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END tie[160]
  PIN tie[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END tie[161]
  PIN tie[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END tie[162]
  PIN tie[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END tie[163]
  PIN tie[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END tie[164]
  PIN tie[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END tie[165]
  PIN tie[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END tie[166]
  PIN tie[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END tie[167]
  PIN tie[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 426.400 4.000 427.000 ;
    END
  END tie[168]
  PIN tie[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END tie[169]
  PIN tie[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END tie[16]
  PIN tie[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END tie[17]
  PIN tie[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END tie[18]
  PIN tie[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END tie[19]
  PIN tie[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END tie[1]
  PIN tie[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END tie[20]
  PIN tie[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END tie[21]
  PIN tie[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END tie[22]
  PIN tie[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END tie[23]
  PIN tie[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END tie[24]
  PIN tie[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END tie[25]
  PIN tie[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END tie[26]
  PIN tie[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END tie[27]
  PIN tie[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END tie[28]
  PIN tie[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END tie[29]
  PIN tie[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END tie[2]
  PIN tie[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END tie[30]
  PIN tie[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END tie[31]
  PIN tie[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END tie[32]
  PIN tie[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END tie[33]
  PIN tie[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END tie[34]
  PIN tie[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END tie[35]
  PIN tie[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END tie[36]
  PIN tie[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END tie[37]
  PIN tie[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END tie[38]
  PIN tie[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END tie[39]
  PIN tie[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END tie[3]
  PIN tie[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END tie[40]
  PIN tie[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END tie[41]
  PIN tie[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END tie[42]
  PIN tie[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END tie[43]
  PIN tie[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END tie[44]
  PIN tie[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END tie[45]
  PIN tie[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END tie[46]
  PIN tie[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END tie[47]
  PIN tie[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END tie[48]
  PIN tie[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END tie[49]
  PIN tie[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END tie[4]
  PIN tie[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END tie[50]
  PIN tie[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END tie[51]
  PIN tie[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END tie[52]
  PIN tie[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END tie[53]
  PIN tie[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END tie[54]
  PIN tie[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END tie[55]
  PIN tie[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END tie[56]
  PIN tie[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END tie[57]
  PIN tie[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END tie[58]
  PIN tie[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END tie[59]
  PIN tie[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END tie[5]
  PIN tie[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END tie[60]
  PIN tie[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END tie[61]
  PIN tie[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END tie[62]
  PIN tie[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END tie[63]
  PIN tie[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END tie[64]
  PIN tie[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END tie[65]
  PIN tie[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END tie[66]
  PIN tie[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END tie[67]
  PIN tie[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END tie[68]
  PIN tie[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END tie[69]
  PIN tie[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END tie[6]
  PIN tie[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END tie[70]
  PIN tie[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END tie[71]
  PIN tie[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END tie[72]
  PIN tie[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END tie[73]
  PIN tie[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END tie[74]
  PIN tie[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END tie[75]
  PIN tie[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END tie[76]
  PIN tie[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END tie[77]
  PIN tie[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END tie[78]
  PIN tie[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END tie[79]
  PIN tie[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END tie[7]
  PIN tie[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END tie[80]
  PIN tie[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END tie[81]
  PIN tie[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END tie[82]
  PIN tie[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END tie[83]
  PIN tie[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END tie[84]
  PIN tie[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END tie[85]
  PIN tie[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END tie[86]
  PIN tie[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END tie[87]
  PIN tie[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END tie[88]
  PIN tie[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END tie[89]
  PIN tie[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END tie[8]
  PIN tie[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END tie[90]
  PIN tie[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END tie[91]
  PIN tie[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END tie[92]
  PIN tie[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END tie[93]
  PIN tie[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END tie[94]
  PIN tie[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END tie[95]
  PIN tie[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 20.440 400.000 21.040 ;
    END
  END tie[96]
  PIN tie[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 61.240 400.000 61.840 ;
    END
  END tie[97]
  PIN tie[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 102.040 400.000 102.640 ;
    END
  END tie[98]
  PIN tie[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 142.840 400.000 143.440 ;
    END
  END tie[99]
  PIN tie[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END tie[9]
  PIN tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 47.640 400.000 48.240 ;
    END
  END tms
  PIN trst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 129.240 400.000 129.840 ;
    END
  END trst
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 438.160 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 438.160 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 438.160 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 438.160 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 438.160 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.995 438.005 ;
      LAYER met1 ;
        RECT 0.990 6.840 399.210 438.160 ;
      LAYER met2 ;
        RECT 1.020 445.720 10.850 446.000 ;
        RECT 11.690 445.720 32.930 446.000 ;
        RECT 33.770 445.720 55.010 446.000 ;
        RECT 55.850 445.720 77.550 446.000 ;
        RECT 78.390 445.720 99.630 446.000 ;
        RECT 100.470 445.720 121.710 446.000 ;
        RECT 122.550 445.720 144.250 446.000 ;
        RECT 145.090 445.720 166.330 446.000 ;
        RECT 167.170 445.720 188.410 446.000 ;
        RECT 189.250 445.720 210.950 446.000 ;
        RECT 211.790 445.720 233.030 446.000 ;
        RECT 233.870 445.720 255.110 446.000 ;
        RECT 255.950 445.720 277.650 446.000 ;
        RECT 278.490 445.720 299.730 446.000 ;
        RECT 300.570 445.720 321.810 446.000 ;
        RECT 322.650 445.720 344.350 446.000 ;
        RECT 345.190 445.720 366.430 446.000 ;
        RECT 367.270 445.720 388.510 446.000 ;
        RECT 389.350 445.720 399.180 446.000 ;
        RECT 1.020 4.280 399.180 445.720 ;
        RECT 1.570 4.000 2.570 4.280 ;
        RECT 3.410 4.000 4.410 4.280 ;
        RECT 5.250 4.000 6.710 4.280 ;
        RECT 7.550 4.000 8.550 4.280 ;
        RECT 9.390 4.000 10.850 4.280 ;
        RECT 11.690 4.000 12.690 4.280 ;
        RECT 13.530 4.000 14.530 4.280 ;
        RECT 15.370 4.000 16.830 4.280 ;
        RECT 17.670 4.000 18.670 4.280 ;
        RECT 19.510 4.000 20.970 4.280 ;
        RECT 21.810 4.000 22.810 4.280 ;
        RECT 23.650 4.000 24.650 4.280 ;
        RECT 25.490 4.000 26.950 4.280 ;
        RECT 27.790 4.000 28.790 4.280 ;
        RECT 29.630 4.000 31.090 4.280 ;
        RECT 31.930 4.000 32.930 4.280 ;
        RECT 33.770 4.000 35.230 4.280 ;
        RECT 36.070 4.000 37.070 4.280 ;
        RECT 37.910 4.000 38.910 4.280 ;
        RECT 39.750 4.000 41.210 4.280 ;
        RECT 42.050 4.000 43.050 4.280 ;
        RECT 43.890 4.000 45.350 4.280 ;
        RECT 46.190 4.000 47.190 4.280 ;
        RECT 48.030 4.000 49.030 4.280 ;
        RECT 49.870 4.000 51.330 4.280 ;
        RECT 52.170 4.000 53.170 4.280 ;
        RECT 54.010 4.000 55.470 4.280 ;
        RECT 56.310 4.000 57.310 4.280 ;
        RECT 58.150 4.000 59.610 4.280 ;
        RECT 60.450 4.000 61.450 4.280 ;
        RECT 62.290 4.000 63.290 4.280 ;
        RECT 64.130 4.000 65.590 4.280 ;
        RECT 66.430 4.000 67.430 4.280 ;
        RECT 68.270 4.000 69.730 4.280 ;
        RECT 70.570 4.000 71.570 4.280 ;
        RECT 72.410 4.000 73.410 4.280 ;
        RECT 74.250 4.000 75.710 4.280 ;
        RECT 76.550 4.000 77.550 4.280 ;
        RECT 78.390 4.000 79.850 4.280 ;
        RECT 80.690 4.000 81.690 4.280 ;
        RECT 82.530 4.000 83.990 4.280 ;
        RECT 84.830 4.000 85.830 4.280 ;
        RECT 86.670 4.000 87.670 4.280 ;
        RECT 88.510 4.000 89.970 4.280 ;
        RECT 90.810 4.000 91.810 4.280 ;
        RECT 92.650 4.000 94.110 4.280 ;
        RECT 94.950 4.000 95.950 4.280 ;
        RECT 96.790 4.000 97.790 4.280 ;
        RECT 98.630 4.000 100.090 4.280 ;
        RECT 100.930 4.000 101.930 4.280 ;
        RECT 102.770 4.000 104.230 4.280 ;
        RECT 105.070 4.000 106.070 4.280 ;
        RECT 106.910 4.000 108.370 4.280 ;
        RECT 109.210 4.000 110.210 4.280 ;
        RECT 111.050 4.000 112.050 4.280 ;
        RECT 112.890 4.000 114.350 4.280 ;
        RECT 115.190 4.000 116.190 4.280 ;
        RECT 117.030 4.000 118.490 4.280 ;
        RECT 119.330 4.000 120.330 4.280 ;
        RECT 121.170 4.000 122.170 4.280 ;
        RECT 123.010 4.000 124.470 4.280 ;
        RECT 125.310 4.000 126.310 4.280 ;
        RECT 127.150 4.000 128.610 4.280 ;
        RECT 129.450 4.000 130.450 4.280 ;
        RECT 131.290 4.000 132.750 4.280 ;
        RECT 133.590 4.000 134.590 4.280 ;
        RECT 135.430 4.000 136.430 4.280 ;
        RECT 137.270 4.000 138.730 4.280 ;
        RECT 139.570 4.000 140.570 4.280 ;
        RECT 141.410 4.000 142.870 4.280 ;
        RECT 143.710 4.000 144.710 4.280 ;
        RECT 145.550 4.000 146.550 4.280 ;
        RECT 147.390 4.000 148.850 4.280 ;
        RECT 149.690 4.000 150.690 4.280 ;
        RECT 151.530 4.000 152.990 4.280 ;
        RECT 153.830 4.000 154.830 4.280 ;
        RECT 155.670 4.000 157.130 4.280 ;
        RECT 157.970 4.000 158.970 4.280 ;
        RECT 159.810 4.000 160.810 4.280 ;
        RECT 161.650 4.000 163.110 4.280 ;
        RECT 163.950 4.000 164.950 4.280 ;
        RECT 165.790 4.000 167.250 4.280 ;
        RECT 168.090 4.000 169.090 4.280 ;
        RECT 169.930 4.000 170.930 4.280 ;
        RECT 171.770 4.000 173.230 4.280 ;
        RECT 174.070 4.000 175.070 4.280 ;
        RECT 175.910 4.000 177.370 4.280 ;
        RECT 178.210 4.000 179.210 4.280 ;
        RECT 180.050 4.000 181.510 4.280 ;
        RECT 182.350 4.000 183.350 4.280 ;
        RECT 184.190 4.000 185.190 4.280 ;
        RECT 186.030 4.000 187.490 4.280 ;
        RECT 188.330 4.000 189.330 4.280 ;
        RECT 190.170 4.000 191.630 4.280 ;
        RECT 192.470 4.000 193.470 4.280 ;
        RECT 194.310 4.000 195.310 4.280 ;
        RECT 196.150 4.000 197.610 4.280 ;
        RECT 198.450 4.000 199.450 4.280 ;
        RECT 200.290 4.000 201.750 4.280 ;
        RECT 202.590 4.000 203.590 4.280 ;
        RECT 204.430 4.000 205.890 4.280 ;
        RECT 206.730 4.000 207.730 4.280 ;
        RECT 208.570 4.000 209.570 4.280 ;
        RECT 210.410 4.000 211.870 4.280 ;
        RECT 212.710 4.000 213.710 4.280 ;
        RECT 214.550 4.000 216.010 4.280 ;
        RECT 216.850 4.000 217.850 4.280 ;
        RECT 218.690 4.000 219.690 4.280 ;
        RECT 220.530 4.000 221.990 4.280 ;
        RECT 222.830 4.000 223.830 4.280 ;
        RECT 224.670 4.000 226.130 4.280 ;
        RECT 226.970 4.000 227.970 4.280 ;
        RECT 228.810 4.000 230.270 4.280 ;
        RECT 231.110 4.000 232.110 4.280 ;
        RECT 232.950 4.000 233.950 4.280 ;
        RECT 234.790 4.000 236.250 4.280 ;
        RECT 237.090 4.000 238.090 4.280 ;
        RECT 238.930 4.000 240.390 4.280 ;
        RECT 241.230 4.000 242.230 4.280 ;
        RECT 243.070 4.000 244.070 4.280 ;
        RECT 244.910 4.000 246.370 4.280 ;
        RECT 247.210 4.000 248.210 4.280 ;
        RECT 249.050 4.000 250.510 4.280 ;
        RECT 251.350 4.000 252.350 4.280 ;
        RECT 253.190 4.000 254.650 4.280 ;
        RECT 255.490 4.000 256.490 4.280 ;
        RECT 257.330 4.000 258.330 4.280 ;
        RECT 259.170 4.000 260.630 4.280 ;
        RECT 261.470 4.000 262.470 4.280 ;
        RECT 263.310 4.000 264.770 4.280 ;
        RECT 265.610 4.000 266.610 4.280 ;
        RECT 267.450 4.000 268.450 4.280 ;
        RECT 269.290 4.000 270.750 4.280 ;
        RECT 271.590 4.000 272.590 4.280 ;
        RECT 273.430 4.000 274.890 4.280 ;
        RECT 275.730 4.000 276.730 4.280 ;
        RECT 277.570 4.000 279.030 4.280 ;
        RECT 279.870 4.000 280.870 4.280 ;
        RECT 281.710 4.000 282.710 4.280 ;
        RECT 283.550 4.000 285.010 4.280 ;
        RECT 285.850 4.000 286.850 4.280 ;
        RECT 287.690 4.000 289.150 4.280 ;
        RECT 289.990 4.000 290.990 4.280 ;
        RECT 291.830 4.000 292.830 4.280 ;
        RECT 293.670 4.000 295.130 4.280 ;
        RECT 295.970 4.000 296.970 4.280 ;
        RECT 297.810 4.000 299.270 4.280 ;
        RECT 300.110 4.000 301.110 4.280 ;
        RECT 301.950 4.000 303.410 4.280 ;
        RECT 304.250 4.000 305.250 4.280 ;
        RECT 306.090 4.000 307.090 4.280 ;
        RECT 307.930 4.000 309.390 4.280 ;
        RECT 310.230 4.000 311.230 4.280 ;
        RECT 312.070 4.000 313.530 4.280 ;
        RECT 314.370 4.000 315.370 4.280 ;
        RECT 316.210 4.000 317.210 4.280 ;
        RECT 318.050 4.000 319.510 4.280 ;
        RECT 320.350 4.000 321.350 4.280 ;
        RECT 322.190 4.000 323.650 4.280 ;
        RECT 324.490 4.000 325.490 4.280 ;
        RECT 326.330 4.000 327.790 4.280 ;
        RECT 328.630 4.000 329.630 4.280 ;
        RECT 330.470 4.000 331.470 4.280 ;
        RECT 332.310 4.000 333.770 4.280 ;
        RECT 334.610 4.000 335.610 4.280 ;
        RECT 336.450 4.000 337.910 4.280 ;
        RECT 338.750 4.000 339.750 4.280 ;
        RECT 340.590 4.000 341.590 4.280 ;
        RECT 342.430 4.000 343.890 4.280 ;
        RECT 344.730 4.000 345.730 4.280 ;
        RECT 346.570 4.000 348.030 4.280 ;
        RECT 348.870 4.000 349.870 4.280 ;
        RECT 350.710 4.000 352.170 4.280 ;
        RECT 353.010 4.000 354.010 4.280 ;
        RECT 354.850 4.000 355.850 4.280 ;
        RECT 356.690 4.000 358.150 4.280 ;
        RECT 358.990 4.000 359.990 4.280 ;
        RECT 360.830 4.000 362.290 4.280 ;
        RECT 363.130 4.000 364.130 4.280 ;
        RECT 364.970 4.000 365.970 4.280 ;
        RECT 366.810 4.000 368.270 4.280 ;
        RECT 369.110 4.000 370.110 4.280 ;
        RECT 370.950 4.000 372.410 4.280 ;
        RECT 373.250 4.000 374.250 4.280 ;
        RECT 375.090 4.000 376.550 4.280 ;
        RECT 377.390 4.000 378.390 4.280 ;
        RECT 379.230 4.000 380.230 4.280 ;
        RECT 381.070 4.000 382.530 4.280 ;
        RECT 383.370 4.000 384.370 4.280 ;
        RECT 385.210 4.000 386.670 4.280 ;
        RECT 387.510 4.000 388.510 4.280 ;
        RECT 389.350 4.000 390.350 4.280 ;
        RECT 391.190 4.000 392.650 4.280 ;
        RECT 393.490 4.000 394.490 4.280 ;
        RECT 395.330 4.000 396.790 4.280 ;
        RECT 397.630 4.000 398.630 4.280 ;
      LAYER met3 ;
        RECT 4.000 443.040 395.600 443.185 ;
        RECT 4.400 442.320 395.600 443.040 ;
        RECT 4.400 441.640 396.000 442.320 ;
        RECT 4.000 430.120 396.000 441.640 ;
        RECT 4.000 428.720 395.600 430.120 ;
        RECT 4.000 427.400 396.000 428.720 ;
        RECT 4.400 426.000 396.000 427.400 ;
        RECT 4.000 416.520 396.000 426.000 ;
        RECT 4.000 415.120 395.600 416.520 ;
        RECT 4.000 411.760 396.000 415.120 ;
        RECT 4.400 410.360 396.000 411.760 ;
        RECT 4.000 402.920 396.000 410.360 ;
        RECT 4.000 401.520 395.600 402.920 ;
        RECT 4.000 396.120 396.000 401.520 ;
        RECT 4.400 394.720 396.000 396.120 ;
        RECT 4.000 389.320 396.000 394.720 ;
        RECT 4.000 387.920 395.600 389.320 ;
        RECT 4.000 380.480 396.000 387.920 ;
        RECT 4.400 379.080 396.000 380.480 ;
        RECT 4.000 375.720 396.000 379.080 ;
        RECT 4.000 374.320 395.600 375.720 ;
        RECT 4.000 365.520 396.000 374.320 ;
        RECT 4.400 364.120 396.000 365.520 ;
        RECT 4.000 362.120 396.000 364.120 ;
        RECT 4.000 360.720 395.600 362.120 ;
        RECT 4.000 349.880 396.000 360.720 ;
        RECT 4.400 348.520 396.000 349.880 ;
        RECT 4.400 348.480 395.600 348.520 ;
        RECT 4.000 347.120 395.600 348.480 ;
        RECT 4.000 334.920 396.000 347.120 ;
        RECT 4.000 334.240 395.600 334.920 ;
        RECT 4.400 333.520 395.600 334.240 ;
        RECT 4.400 332.840 396.000 333.520 ;
        RECT 4.000 321.320 396.000 332.840 ;
        RECT 4.000 319.920 395.600 321.320 ;
        RECT 4.000 318.600 396.000 319.920 ;
        RECT 4.400 317.200 396.000 318.600 ;
        RECT 4.000 307.720 396.000 317.200 ;
        RECT 4.000 306.320 395.600 307.720 ;
        RECT 4.000 302.960 396.000 306.320 ;
        RECT 4.400 301.560 396.000 302.960 ;
        RECT 4.000 294.120 396.000 301.560 ;
        RECT 4.000 292.720 395.600 294.120 ;
        RECT 4.000 287.320 396.000 292.720 ;
        RECT 4.400 285.920 396.000 287.320 ;
        RECT 4.000 280.520 396.000 285.920 ;
        RECT 4.000 279.120 395.600 280.520 ;
        RECT 4.000 272.360 396.000 279.120 ;
        RECT 4.400 270.960 396.000 272.360 ;
        RECT 4.000 266.920 396.000 270.960 ;
        RECT 4.000 265.520 395.600 266.920 ;
        RECT 4.000 256.720 396.000 265.520 ;
        RECT 4.400 255.320 396.000 256.720 ;
        RECT 4.000 253.320 396.000 255.320 ;
        RECT 4.000 251.920 395.600 253.320 ;
        RECT 4.000 241.080 396.000 251.920 ;
        RECT 4.400 239.720 396.000 241.080 ;
        RECT 4.400 239.680 395.600 239.720 ;
        RECT 4.000 238.320 395.600 239.680 ;
        RECT 4.000 225.440 396.000 238.320 ;
        RECT 4.400 224.040 395.600 225.440 ;
        RECT 4.000 211.840 396.000 224.040 ;
        RECT 4.000 210.440 395.600 211.840 ;
        RECT 4.000 209.800 396.000 210.440 ;
        RECT 4.400 208.400 396.000 209.800 ;
        RECT 4.000 198.240 396.000 208.400 ;
        RECT 4.000 196.840 395.600 198.240 ;
        RECT 4.000 194.160 396.000 196.840 ;
        RECT 4.400 192.760 396.000 194.160 ;
        RECT 4.000 184.640 396.000 192.760 ;
        RECT 4.000 183.240 395.600 184.640 ;
        RECT 4.000 179.200 396.000 183.240 ;
        RECT 4.400 177.800 396.000 179.200 ;
        RECT 4.000 171.040 396.000 177.800 ;
        RECT 4.000 169.640 395.600 171.040 ;
        RECT 4.000 163.560 396.000 169.640 ;
        RECT 4.400 162.160 396.000 163.560 ;
        RECT 4.000 157.440 396.000 162.160 ;
        RECT 4.000 156.040 395.600 157.440 ;
        RECT 4.000 147.920 396.000 156.040 ;
        RECT 4.400 146.520 396.000 147.920 ;
        RECT 4.000 143.840 396.000 146.520 ;
        RECT 4.000 142.440 395.600 143.840 ;
        RECT 4.000 132.280 396.000 142.440 ;
        RECT 4.400 130.880 396.000 132.280 ;
        RECT 4.000 130.240 396.000 130.880 ;
        RECT 4.000 128.840 395.600 130.240 ;
        RECT 4.000 116.640 396.000 128.840 ;
        RECT 4.400 115.240 395.600 116.640 ;
        RECT 4.000 103.040 396.000 115.240 ;
        RECT 4.000 101.640 395.600 103.040 ;
        RECT 4.000 101.000 396.000 101.640 ;
        RECT 4.400 99.600 396.000 101.000 ;
        RECT 4.000 89.440 396.000 99.600 ;
        RECT 4.000 88.040 395.600 89.440 ;
        RECT 4.000 86.040 396.000 88.040 ;
        RECT 4.400 84.640 396.000 86.040 ;
        RECT 4.000 75.840 396.000 84.640 ;
        RECT 4.000 74.440 395.600 75.840 ;
        RECT 4.000 70.400 396.000 74.440 ;
        RECT 4.400 69.000 396.000 70.400 ;
        RECT 4.000 62.240 396.000 69.000 ;
        RECT 4.000 60.840 395.600 62.240 ;
        RECT 4.000 54.760 396.000 60.840 ;
        RECT 4.400 53.360 396.000 54.760 ;
        RECT 4.000 48.640 396.000 53.360 ;
        RECT 4.000 47.240 395.600 48.640 ;
        RECT 4.000 39.120 396.000 47.240 ;
        RECT 4.400 37.720 396.000 39.120 ;
        RECT 4.000 35.040 396.000 37.720 ;
        RECT 4.000 33.640 395.600 35.040 ;
        RECT 4.000 23.480 396.000 33.640 ;
        RECT 4.400 22.080 396.000 23.480 ;
        RECT 4.000 21.440 396.000 22.080 ;
        RECT 4.000 20.040 395.600 21.440 ;
        RECT 4.000 8.520 396.000 20.040 ;
        RECT 4.400 7.840 396.000 8.520 ;
        RECT 4.400 7.120 395.600 7.840 ;
        RECT 4.000 6.975 395.600 7.120 ;
  END
END user_proj_top
END LIBRARY

