magic
tech sky130A
magscale 1 2
timestamp 1612285914
<< obsli1 >>
rect 1104 2159 78999 87601
<< obsm1 >>
rect 198 1368 79842 87632
<< metal2 >>
rect 2226 89200 2282 90000
rect 6642 89200 6698 90000
rect 11058 89200 11114 90000
rect 15566 89200 15622 90000
rect 19982 89200 20038 90000
rect 24398 89200 24454 90000
rect 28906 89200 28962 90000
rect 33322 89200 33378 90000
rect 37738 89200 37794 90000
rect 42246 89200 42302 90000
rect 46662 89200 46718 90000
rect 51078 89200 51134 90000
rect 55586 89200 55642 90000
rect 60002 89200 60058 90000
rect 64418 89200 64474 90000
rect 68926 89200 68982 90000
rect 73342 89200 73398 90000
rect 77758 89200 77814 90000
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20902 0 20958 800
rect 21270 0 21326 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22926 0 22982 800
rect 23294 0 23350 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24950 0 25006 800
rect 25318 0 25374 800
rect 25778 0 25834 800
rect 26146 0 26202 800
rect 26606 0 26662 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29826 0 29882 800
rect 30194 0 30250 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32678 0 32734 800
rect 33046 0 33102 800
rect 33506 0 33562 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34702 0 34758 800
rect 35070 0 35126 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36726 0 36782 800
rect 37094 0 37150 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38382 0 38438 800
rect 38750 0 38806 800
rect 39118 0 39174 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41234 0 41290 800
rect 41602 0 41658 800
rect 41970 0 42026 800
rect 42430 0 42486 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43994 0 44050 800
rect 44454 0 44510 800
rect 44822 0 44878 800
rect 45282 0 45338 800
rect 45650 0 45706 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46846 0 46902 800
rect 47306 0 47362 800
rect 47674 0 47730 800
rect 48134 0 48190 800
rect 48502 0 48558 800
rect 48870 0 48926 800
rect 49330 0 49386 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 50526 0 50582 800
rect 50986 0 51042 800
rect 51354 0 51410 800
rect 51722 0 51778 800
rect 52182 0 52238 800
rect 52550 0 52606 800
rect 53010 0 53066 800
rect 53378 0 53434 800
rect 53746 0 53802 800
rect 54206 0 54262 800
rect 54574 0 54630 800
rect 55034 0 55090 800
rect 55402 0 55458 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56598 0 56654 800
rect 57058 0 57114 800
rect 57426 0 57482 800
rect 57886 0 57942 800
rect 58254 0 58310 800
rect 58622 0 58678 800
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59910 0 59966 800
rect 60278 0 60334 800
rect 60738 0 60794 800
rect 61106 0 61162 800
rect 61474 0 61530 800
rect 61934 0 61990 800
rect 62302 0 62358 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63958 0 64014 800
rect 64326 0 64382 800
rect 64786 0 64842 800
rect 65154 0 65210 800
rect 65614 0 65670 800
rect 65982 0 66038 800
rect 66350 0 66406 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68374 0 68430 800
rect 68834 0 68890 800
rect 69202 0 69258 800
rect 69662 0 69718 800
rect 70030 0 70086 800
rect 70490 0 70546 800
rect 70858 0 70914 800
rect 71226 0 71282 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72514 0 72570 800
rect 72882 0 72938 800
rect 73250 0 73306 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75366 0 75422 800
rect 75734 0 75790 800
rect 76102 0 76158 800
rect 76562 0 76618 800
rect 76930 0 76986 800
rect 77390 0 77446 800
rect 77758 0 77814 800
rect 78126 0 78182 800
rect 78586 0 78642 800
rect 78954 0 79010 800
rect 79414 0 79470 800
rect 79782 0 79838 800
<< obsm2 >>
rect 204 89144 2170 89200
rect 2338 89144 6586 89200
rect 6754 89144 11002 89200
rect 11170 89144 15510 89200
rect 15678 89144 19926 89200
rect 20094 89144 24342 89200
rect 24510 89144 28850 89200
rect 29018 89144 33266 89200
rect 33434 89144 37682 89200
rect 37850 89144 42190 89200
rect 42358 89144 46606 89200
rect 46774 89144 51022 89200
rect 51190 89144 55530 89200
rect 55698 89144 59946 89200
rect 60114 89144 64362 89200
rect 64530 89144 68870 89200
rect 69038 89144 73286 89200
rect 73454 89144 77702 89200
rect 77870 89144 79836 89200
rect 204 856 79836 89144
rect 314 800 514 856
rect 682 800 882 856
rect 1050 800 1342 856
rect 1510 800 1710 856
rect 1878 800 2170 856
rect 2338 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3366 856
rect 3534 800 3734 856
rect 3902 800 4194 856
rect 4362 800 4562 856
rect 4730 800 4930 856
rect 5098 800 5390 856
rect 5558 800 5758 856
rect 5926 800 6218 856
rect 6386 800 6586 856
rect 6754 800 7046 856
rect 7214 800 7414 856
rect 7582 800 7782 856
rect 7950 800 8242 856
rect 8410 800 8610 856
rect 8778 800 9070 856
rect 9238 800 9438 856
rect 9606 800 9806 856
rect 9974 800 10266 856
rect 10434 800 10634 856
rect 10802 800 11094 856
rect 11262 800 11462 856
rect 11630 800 11922 856
rect 12090 800 12290 856
rect 12458 800 12658 856
rect 12826 800 13118 856
rect 13286 800 13486 856
rect 13654 800 13946 856
rect 14114 800 14314 856
rect 14482 800 14682 856
rect 14850 800 15142 856
rect 15310 800 15510 856
rect 15678 800 15970 856
rect 16138 800 16338 856
rect 16506 800 16798 856
rect 16966 800 17166 856
rect 17334 800 17534 856
rect 17702 800 17994 856
rect 18162 800 18362 856
rect 18530 800 18822 856
rect 18990 800 19190 856
rect 19358 800 19558 856
rect 19726 800 20018 856
rect 20186 800 20386 856
rect 20554 800 20846 856
rect 21014 800 21214 856
rect 21382 800 21674 856
rect 21842 800 22042 856
rect 22210 800 22410 856
rect 22578 800 22870 856
rect 23038 800 23238 856
rect 23406 800 23698 856
rect 23866 800 24066 856
rect 24234 800 24434 856
rect 24602 800 24894 856
rect 25062 800 25262 856
rect 25430 800 25722 856
rect 25890 800 26090 856
rect 26258 800 26550 856
rect 26718 800 26918 856
rect 27086 800 27286 856
rect 27454 800 27746 856
rect 27914 800 28114 856
rect 28282 800 28574 856
rect 28742 800 28942 856
rect 29110 800 29310 856
rect 29478 800 29770 856
rect 29938 800 30138 856
rect 30306 800 30598 856
rect 30766 800 30966 856
rect 31134 800 31426 856
rect 31594 800 31794 856
rect 31962 800 32162 856
rect 32330 800 32622 856
rect 32790 800 32990 856
rect 33158 800 33450 856
rect 33618 800 33818 856
rect 33986 800 34186 856
rect 34354 800 34646 856
rect 34814 800 35014 856
rect 35182 800 35474 856
rect 35642 800 35842 856
rect 36010 800 36302 856
rect 36470 800 36670 856
rect 36838 800 37038 856
rect 37206 800 37498 856
rect 37666 800 37866 856
rect 38034 800 38326 856
rect 38494 800 38694 856
rect 38862 800 39062 856
rect 39230 800 39522 856
rect 39690 800 39890 856
rect 40058 800 40350 856
rect 40518 800 40718 856
rect 40886 800 41178 856
rect 41346 800 41546 856
rect 41714 800 41914 856
rect 42082 800 42374 856
rect 42542 800 42742 856
rect 42910 800 43202 856
rect 43370 800 43570 856
rect 43738 800 43938 856
rect 44106 800 44398 856
rect 44566 800 44766 856
rect 44934 800 45226 856
rect 45394 800 45594 856
rect 45762 800 46054 856
rect 46222 800 46422 856
rect 46590 800 46790 856
rect 46958 800 47250 856
rect 47418 800 47618 856
rect 47786 800 48078 856
rect 48246 800 48446 856
rect 48614 800 48814 856
rect 48982 800 49274 856
rect 49442 800 49642 856
rect 49810 800 50102 856
rect 50270 800 50470 856
rect 50638 800 50930 856
rect 51098 800 51298 856
rect 51466 800 51666 856
rect 51834 800 52126 856
rect 52294 800 52494 856
rect 52662 800 52954 856
rect 53122 800 53322 856
rect 53490 800 53690 856
rect 53858 800 54150 856
rect 54318 800 54518 856
rect 54686 800 54978 856
rect 55146 800 55346 856
rect 55514 800 55806 856
rect 55974 800 56174 856
rect 56342 800 56542 856
rect 56710 800 57002 856
rect 57170 800 57370 856
rect 57538 800 57830 856
rect 57998 800 58198 856
rect 58366 800 58566 856
rect 58734 800 59026 856
rect 59194 800 59394 856
rect 59562 800 59854 856
rect 60022 800 60222 856
rect 60390 800 60682 856
rect 60850 800 61050 856
rect 61218 800 61418 856
rect 61586 800 61878 856
rect 62046 800 62246 856
rect 62414 800 62706 856
rect 62874 800 63074 856
rect 63242 800 63442 856
rect 63610 800 63902 856
rect 64070 800 64270 856
rect 64438 800 64730 856
rect 64898 800 65098 856
rect 65266 800 65558 856
rect 65726 800 65926 856
rect 66094 800 66294 856
rect 66462 800 66754 856
rect 66922 800 67122 856
rect 67290 800 67582 856
rect 67750 800 67950 856
rect 68118 800 68318 856
rect 68486 800 68778 856
rect 68946 800 69146 856
rect 69314 800 69606 856
rect 69774 800 69974 856
rect 70142 800 70434 856
rect 70602 800 70802 856
rect 70970 800 71170 856
rect 71338 800 71630 856
rect 71798 800 71998 856
rect 72166 800 72458 856
rect 72626 800 72826 856
rect 72994 800 73194 856
rect 73362 800 73654 856
rect 73822 800 74022 856
rect 74190 800 74482 856
rect 74650 800 74850 856
rect 75018 800 75310 856
rect 75478 800 75678 856
rect 75846 800 76046 856
rect 76214 800 76506 856
rect 76674 800 76874 856
rect 77042 800 77334 856
rect 77502 800 77702 856
rect 77870 800 78070 856
rect 78238 800 78530 856
rect 78698 800 78898 856
rect 79066 800 79358 856
rect 79526 800 79726 856
<< metal3 >>
rect 0 88408 800 88528
rect 79200 88544 80000 88664
rect 79200 85824 80000 85944
rect 0 85280 800 85400
rect 79200 83104 80000 83224
rect 0 82152 800 82272
rect 79200 80384 80000 80504
rect 0 79024 800 79144
rect 79200 77664 80000 77784
rect 0 75896 800 76016
rect 79200 74944 80000 75064
rect 0 72904 800 73024
rect 79200 72224 80000 72344
rect 0 69776 800 69896
rect 79200 69504 80000 69624
rect 0 66648 800 66768
rect 79200 66784 80000 66904
rect 79200 64064 80000 64184
rect 0 63520 800 63640
rect 79200 61344 80000 61464
rect 0 60392 800 60512
rect 79200 58624 80000 58744
rect 0 57264 800 57384
rect 79200 55904 80000 56024
rect 0 54272 800 54392
rect 79200 53184 80000 53304
rect 0 51144 800 51264
rect 79200 50464 80000 50584
rect 0 48016 800 48136
rect 79200 47744 80000 47864
rect 0 44888 800 45008
rect 79200 44888 80000 45008
rect 79200 42168 80000 42288
rect 0 41760 800 41880
rect 79200 39448 80000 39568
rect 0 38632 800 38752
rect 79200 36728 80000 36848
rect 0 35640 800 35760
rect 79200 34008 80000 34128
rect 0 32512 800 32632
rect 79200 31288 80000 31408
rect 0 29384 800 29504
rect 79200 28568 80000 28688
rect 0 26256 800 26376
rect 79200 25848 80000 25968
rect 0 23128 800 23248
rect 79200 23128 80000 23248
rect 79200 20408 80000 20528
rect 0 20000 800 20120
rect 79200 17688 80000 17808
rect 0 17008 800 17128
rect 79200 14968 80000 15088
rect 0 13880 800 14000
rect 79200 12248 80000 12368
rect 0 10752 800 10872
rect 79200 9528 80000 9648
rect 0 7624 800 7744
rect 79200 6808 80000 6928
rect 0 4496 800 4616
rect 79200 4088 80000 4208
rect 0 1504 800 1624
rect 79200 1368 80000 1488
<< obsm3 >>
rect 800 88608 79120 88637
rect 880 88464 79120 88608
rect 880 88328 79200 88464
rect 800 86024 79200 88328
rect 800 85744 79120 86024
rect 800 85480 79200 85744
rect 880 85200 79200 85480
rect 800 83304 79200 85200
rect 800 83024 79120 83304
rect 800 82352 79200 83024
rect 880 82072 79200 82352
rect 800 80584 79200 82072
rect 800 80304 79120 80584
rect 800 79224 79200 80304
rect 880 78944 79200 79224
rect 800 77864 79200 78944
rect 800 77584 79120 77864
rect 800 76096 79200 77584
rect 880 75816 79200 76096
rect 800 75144 79200 75816
rect 800 74864 79120 75144
rect 800 73104 79200 74864
rect 880 72824 79200 73104
rect 800 72424 79200 72824
rect 800 72144 79120 72424
rect 800 69976 79200 72144
rect 880 69704 79200 69976
rect 880 69696 79120 69704
rect 800 69424 79120 69696
rect 800 66984 79200 69424
rect 800 66848 79120 66984
rect 880 66704 79120 66848
rect 880 66568 79200 66704
rect 800 64264 79200 66568
rect 800 63984 79120 64264
rect 800 63720 79200 63984
rect 880 63440 79200 63720
rect 800 61544 79200 63440
rect 800 61264 79120 61544
rect 800 60592 79200 61264
rect 880 60312 79200 60592
rect 800 58824 79200 60312
rect 800 58544 79120 58824
rect 800 57464 79200 58544
rect 880 57184 79200 57464
rect 800 56104 79200 57184
rect 800 55824 79120 56104
rect 800 54472 79200 55824
rect 880 54192 79200 54472
rect 800 53384 79200 54192
rect 800 53104 79120 53384
rect 800 51344 79200 53104
rect 880 51064 79200 51344
rect 800 50664 79200 51064
rect 800 50384 79120 50664
rect 800 48216 79200 50384
rect 880 47944 79200 48216
rect 880 47936 79120 47944
rect 800 47664 79120 47936
rect 800 45088 79200 47664
rect 880 44808 79120 45088
rect 800 42368 79200 44808
rect 800 42088 79120 42368
rect 800 41960 79200 42088
rect 880 41680 79200 41960
rect 800 39648 79200 41680
rect 800 39368 79120 39648
rect 800 38832 79200 39368
rect 880 38552 79200 38832
rect 800 36928 79200 38552
rect 800 36648 79120 36928
rect 800 35840 79200 36648
rect 880 35560 79200 35840
rect 800 34208 79200 35560
rect 800 33928 79120 34208
rect 800 32712 79200 33928
rect 880 32432 79200 32712
rect 800 31488 79200 32432
rect 800 31208 79120 31488
rect 800 29584 79200 31208
rect 880 29304 79200 29584
rect 800 28768 79200 29304
rect 800 28488 79120 28768
rect 800 26456 79200 28488
rect 880 26176 79200 26456
rect 800 26048 79200 26176
rect 800 25768 79120 26048
rect 800 23328 79200 25768
rect 880 23048 79120 23328
rect 800 20608 79200 23048
rect 800 20328 79120 20608
rect 800 20200 79200 20328
rect 880 19920 79200 20200
rect 800 17888 79200 19920
rect 800 17608 79120 17888
rect 800 17208 79200 17608
rect 880 16928 79200 17208
rect 800 15168 79200 16928
rect 800 14888 79120 15168
rect 800 14080 79200 14888
rect 880 13800 79200 14080
rect 800 12448 79200 13800
rect 800 12168 79120 12448
rect 800 10952 79200 12168
rect 880 10672 79200 10952
rect 800 9728 79200 10672
rect 800 9448 79120 9728
rect 800 7824 79200 9448
rect 880 7544 79200 7824
rect 800 7008 79200 7544
rect 800 6728 79120 7008
rect 800 4696 79200 6728
rect 880 4416 79200 4696
rect 800 4288 79200 4416
rect 800 4008 79120 4288
rect 800 1704 79200 4008
rect 880 1568 79200 1704
rect 880 1424 79120 1568
rect 800 1395 79120 1424
<< metal4 >>
rect 4208 2128 4528 87632
rect 19568 2128 19888 87632
rect 34928 2128 35248 87632
rect 50288 2128 50608 87632
rect 65648 2128 65968 87632
<< labels >>
rlabel metal2 s 202 0 258 800 6 clk
port 1 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 done
port 2 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 mc[0]
port 3 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 mc[10]
port 4 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 mc[11]
port 5 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 mc[12]
port 6 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 mc[13]
port 7 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 mc[14]
port 8 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 mc[15]
port 9 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 mc[16]
port 10 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 mc[17]
port 11 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 mc[18]
port 12 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 mc[19]
port 13 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 mc[1]
port 14 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 mc[20]
port 15 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 mc[21]
port 16 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 mc[22]
port 17 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 mc[23]
port 18 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 mc[24]
port 19 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 mc[25]
port 20 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 mc[26]
port 21 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 mc[27]
port 22 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 mc[28]
port 23 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 mc[29]
port 24 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 mc[2]
port 25 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 mc[30]
port 26 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 mc[31]
port 27 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 mc[3]
port 28 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 mc[4]
port 29 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 mc[5]
port 30 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 mc[6]
port 31 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 mc[7]
port 32 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 mc[8]
port 33 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 mc[9]
port 34 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 mp[0]
port 35 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 mp[10]
port 36 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 mp[11]
port 37 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 mp[12]
port 38 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 mp[13]
port 39 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 mp[14]
port 40 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 mp[15]
port 41 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 mp[16]
port 42 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 mp[17]
port 43 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 mp[18]
port 44 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 mp[19]
port 45 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 mp[1]
port 46 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 mp[20]
port 47 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 mp[21]
port 48 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 mp[22]
port 49 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 mp[23]
port 50 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 mp[24]
port 51 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 mp[25]
port 52 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 mp[26]
port 53 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 mp[27]
port 54 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 mp[28]
port 55 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 mp[29]
port 56 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 mp[2]
port 57 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 mp[30]
port 58 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 mp[31]
port 59 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 mp[3]
port 60 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 mp[4]
port 61 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 mp[5]
port 62 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 mp[6]
port 63 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 mp[7]
port 64 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 mp[8]
port 65 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 mp[9]
port 66 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 prod[0]
port 67 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 prod[10]
port 68 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 prod[11]
port 69 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 prod[12]
port 70 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 prod[13]
port 71 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 prod[14]
port 72 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 prod[15]
port 73 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 prod[16]
port 74 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 prod[17]
port 75 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 prod[18]
port 76 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 prod[19]
port 77 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 prod[1]
port 78 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 prod[20]
port 79 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 prod[21]
port 80 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 prod[22]
port 81 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 prod[23]
port 82 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 prod[24]
port 83 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 prod[25]
port 84 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 prod[26]
port 85 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 prod[27]
port 86 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 prod[28]
port 87 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 prod[29]
port 88 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 prod[2]
port 89 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 prod[30]
port 90 nsew signal output
rlabel metal2 s 79782 0 79838 800 6 prod[31]
port 91 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 prod[3]
port 92 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 prod[4]
port 93 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 prod[5]
port 94 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 prod[6]
port 95 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 prod[7]
port 96 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 prod[8]
port 97 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 prod[9]
port 98 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 prod_sel
port 99 nsew signal input
rlabel metal2 s 570 0 626 800 6 rst
port 100 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 start
port 101 nsew signal input
rlabel metal3 s 79200 1368 80000 1488 6 tck
port 102 nsew signal input
rlabel metal3 s 79200 17688 80000 17808 6 tdi
port 103 nsew signal input
rlabel metal3 s 79200 34008 80000 34128 6 tdo
port 104 nsew signal output
rlabel metal3 s 79200 36728 80000 36848 6 tdo_paden_o
port 105 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 tie[0]
port 106 nsew signal output
rlabel metal3 s 79200 39448 80000 39568 6 tie[100]
port 107 nsew signal output
rlabel metal3 s 79200 42168 80000 42288 6 tie[101]
port 108 nsew signal output
rlabel metal3 s 79200 44888 80000 45008 6 tie[102]
port 109 nsew signal output
rlabel metal3 s 79200 47744 80000 47864 6 tie[103]
port 110 nsew signal output
rlabel metal3 s 79200 50464 80000 50584 6 tie[104]
port 111 nsew signal output
rlabel metal3 s 79200 53184 80000 53304 6 tie[105]
port 112 nsew signal output
rlabel metal3 s 79200 55904 80000 56024 6 tie[106]
port 113 nsew signal output
rlabel metal3 s 79200 58624 80000 58744 6 tie[107]
port 114 nsew signal output
rlabel metal3 s 79200 61344 80000 61464 6 tie[108]
port 115 nsew signal output
rlabel metal3 s 79200 64064 80000 64184 6 tie[109]
port 116 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 tie[10]
port 117 nsew signal output
rlabel metal2 s 2226 89200 2282 90000 6 tie[110]
port 118 nsew signal output
rlabel metal2 s 6642 89200 6698 90000 6 tie[111]
port 119 nsew signal output
rlabel metal2 s 11058 89200 11114 90000 6 tie[112]
port 120 nsew signal output
rlabel metal2 s 15566 89200 15622 90000 6 tie[113]
port 121 nsew signal output
rlabel metal2 s 19982 89200 20038 90000 6 tie[114]
port 122 nsew signal output
rlabel metal2 s 24398 89200 24454 90000 6 tie[115]
port 123 nsew signal output
rlabel metal2 s 28906 89200 28962 90000 6 tie[116]
port 124 nsew signal output
rlabel metal2 s 33322 89200 33378 90000 6 tie[117]
port 125 nsew signal output
rlabel metal2 s 37738 89200 37794 90000 6 tie[118]
port 126 nsew signal output
rlabel metal3 s 0 1504 800 1624 6 tie[119]
port 127 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 tie[11]
port 128 nsew signal output
rlabel metal3 s 0 4496 800 4616 6 tie[120]
port 129 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 tie[121]
port 130 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 tie[122]
port 131 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 tie[123]
port 132 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 tie[124]
port 133 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 tie[125]
port 134 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 tie[126]
port 135 nsew signal output
rlabel metal3 s 0 26256 800 26376 6 tie[127]
port 136 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 tie[128]
port 137 nsew signal output
rlabel metal3 s 0 32512 800 32632 6 tie[129]
port 138 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 tie[12]
port 139 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 tie[130]
port 140 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 tie[131]
port 141 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 tie[132]
port 142 nsew signal output
rlabel metal3 s 79200 6808 80000 6928 6 tie[133]
port 143 nsew signal output
rlabel metal3 s 79200 14968 80000 15088 6 tie[134]
port 144 nsew signal output
rlabel metal3 s 79200 23128 80000 23248 6 tie[135]
port 145 nsew signal output
rlabel metal3 s 79200 31288 80000 31408 6 tie[136]
port 146 nsew signal output
rlabel metal3 s 79200 66784 80000 66904 6 tie[137]
port 147 nsew signal output
rlabel metal3 s 79200 69504 80000 69624 6 tie[138]
port 148 nsew signal output
rlabel metal3 s 79200 72224 80000 72344 6 tie[139]
port 149 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 tie[13]
port 150 nsew signal output
rlabel metal3 s 79200 74944 80000 75064 6 tie[140]
port 151 nsew signal output
rlabel metal3 s 79200 77664 80000 77784 6 tie[141]
port 152 nsew signal output
rlabel metal3 s 79200 80384 80000 80504 6 tie[142]
port 153 nsew signal output
rlabel metal3 s 79200 83104 80000 83224 6 tie[143]
port 154 nsew signal output
rlabel metal3 s 79200 85824 80000 85944 6 tie[144]
port 155 nsew signal output
rlabel metal3 s 79200 88544 80000 88664 6 tie[145]
port 156 nsew signal output
rlabel metal2 s 42246 89200 42302 90000 6 tie[146]
port 157 nsew signal output
rlabel metal2 s 46662 89200 46718 90000 6 tie[147]
port 158 nsew signal output
rlabel metal2 s 51078 89200 51134 90000 6 tie[148]
port 159 nsew signal output
rlabel metal2 s 55586 89200 55642 90000 6 tie[149]
port 160 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 tie[14]
port 161 nsew signal output
rlabel metal2 s 60002 89200 60058 90000 6 tie[150]
port 162 nsew signal output
rlabel metal2 s 64418 89200 64474 90000 6 tie[151]
port 163 nsew signal output
rlabel metal2 s 68926 89200 68982 90000 6 tie[152]
port 164 nsew signal output
rlabel metal2 s 73342 89200 73398 90000 6 tie[153]
port 165 nsew signal output
rlabel metal2 s 77758 89200 77814 90000 6 tie[154]
port 166 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 tie[155]
port 167 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 tie[156]
port 168 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 tie[157]
port 169 nsew signal output
rlabel metal3 s 0 54272 800 54392 6 tie[158]
port 170 nsew signal output
rlabel metal3 s 0 57264 800 57384 6 tie[159]
port 171 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 tie[15]
port 172 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 tie[160]
port 173 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 tie[161]
port 174 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 tie[162]
port 175 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 tie[163]
port 176 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 tie[164]
port 177 nsew signal output
rlabel metal3 s 0 75896 800 76016 6 tie[165]
port 178 nsew signal output
rlabel metal3 s 0 79024 800 79144 6 tie[166]
port 179 nsew signal output
rlabel metal3 s 0 82152 800 82272 6 tie[167]
port 180 nsew signal output
rlabel metal3 s 0 85280 800 85400 6 tie[168]
port 181 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 tie[169]
port 182 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 tie[16]
port 183 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 tie[17]
port 184 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 tie[18]
port 185 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 tie[19]
port 186 nsew signal output
rlabel metal2 s 10690 0 10746 800 6 tie[1]
port 187 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 tie[20]
port 188 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 tie[21]
port 189 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 tie[22]
port 190 nsew signal output
rlabel metal2 s 3422 0 3478 800 6 tie[23]
port 191 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 tie[24]
port 192 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 tie[25]
port 193 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 tie[26]
port 194 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 tie[27]
port 195 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 tie[28]
port 196 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 tie[29]
port 197 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 tie[2]
port 198 nsew signal output
rlabel metal2 s 938 0 994 800 6 tie[30]
port 199 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 tie[31]
port 200 nsew signal output
rlabel metal2 s 1766 0 1822 800 6 tie[32]
port 201 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 tie[33]
port 202 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 tie[34]
port 203 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 tie[35]
port 204 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 tie[36]
port 205 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 tie[37]
port 206 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 tie[38]
port 207 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 tie[39]
port 208 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 tie[3]
port 209 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 tie[40]
port 210 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 tie[41]
port 211 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 tie[42]
port 212 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 tie[43]
port 213 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 tie[44]
port 214 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 tie[45]
port 215 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 tie[46]
port 216 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 tie[47]
port 217 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 tie[48]
port 218 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 tie[49]
port 219 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 tie[4]
port 220 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 tie[50]
port 221 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 tie[51]
port 222 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 tie[52]
port 223 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 tie[53]
port 224 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 tie[54]
port 225 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 tie[55]
port 226 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 tie[56]
port 227 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 tie[57]
port 228 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 tie[58]
port 229 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 tie[59]
port 230 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 tie[5]
port 231 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 tie[60]
port 232 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 tie[61]
port 233 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 tie[62]
port 234 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 tie[63]
port 235 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 tie[64]
port 236 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 tie[65]
port 237 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 tie[66]
port 238 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 tie[67]
port 239 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 tie[68]
port 240 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 tie[69]
port 241 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 tie[6]
port 242 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 tie[70]
port 243 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 tie[71]
port 244 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 tie[72]
port 245 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 tie[73]
port 246 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 tie[74]
port 247 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 tie[75]
port 248 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 tie[76]
port 249 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 tie[77]
port 250 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 tie[78]
port 251 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 tie[79]
port 252 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 tie[7]
port 253 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 tie[80]
port 254 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 tie[81]
port 255 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 tie[82]
port 256 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 tie[83]
port 257 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 tie[84]
port 258 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 tie[85]
port 259 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 tie[86]
port 260 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 tie[87]
port 261 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 tie[88]
port 262 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 tie[89]
port 263 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 tie[8]
port 264 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 tie[90]
port 265 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 tie[91]
port 266 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 tie[92]
port 267 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 tie[93]
port 268 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 tie[94]
port 269 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 tie[95]
port 270 nsew signal output
rlabel metal3 s 79200 4088 80000 4208 6 tie[96]
port 271 nsew signal output
rlabel metal3 s 79200 12248 80000 12368 6 tie[97]
port 272 nsew signal output
rlabel metal3 s 79200 20408 80000 20528 6 tie[98]
port 273 nsew signal output
rlabel metal3 s 79200 28568 80000 28688 6 tie[99]
port 274 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 tie[9]
port 275 nsew signal output
rlabel metal3 s 79200 9528 80000 9648 6 tms
port 276 nsew signal input
rlabel metal3 s 79200 25848 80000 25968 6 trst
port 277 nsew signal input
rlabel metal4 s 65648 2128 65968 87632 6 VPWR
port 278 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 87632 6 VPWR
port 279 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 87632 6 VPWR
port 280 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 87632 6 VGND
port 281 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 87632 6 VGND
port 282 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 80000 90000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_top/runs/user_proj_top/results/magic/user_proj_top.gds
string GDS_END 9293124
string GDS_START 265700
<< end >>

